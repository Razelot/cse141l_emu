// A synchronous instruction memory
`timescale 1ns / 1ps

module instr_mem #(parameter rom_size = 512, parameter instr_width = 9)
(
  input [$clog2(rom_size):0] instr_addr,
  output [instr_width-1:0] instr_out
  );

  // Store instructions in memory
  logic [instr_width-1:0] rom [rom_size-1:0];

  assign instr_out = rom[instr_addr];

  // FOR TESTING
assign rom[0] = 'b001010110;assign rom[1] = 'b001000110;assign rom[2] = 'b111010110;assign rom[3] = 'b001010110;assign rom[4] = 'b111010110;assign rom[5] = 'b001010110;assign rom[6] = 'b111010110;assign rom[7] = 'b001010110;assign rom[8] = 'b111010110;assign rom[9] = 'b001010110;assign rom[10] = 'b111010110;assign rom[11] = 'b001010110;assign rom[12] = 'b111010110;assign rom[13] = 'b001010110;assign rom[14] = 'b111010110;assign rom[15] = 'b001010110;assign rom[16] = 'b101000000;assign rom[17] = 'b001011010;assign rom[18] = 'b001100101;assign rom[19] = 'b001000111;assign rom[20] = 'b001000110;assign rom[21] = 'b001000110;assign rom[22] = 'b001000110;assign rom[23] = 'b001000110;assign rom[24] = 'b001000110;assign rom[25] = 'b001000110;assign rom[26] = 'b001000110;assign rom[27] = 'b001000110;assign rom[28] = 'b001000110;assign rom[29] = 'b001001010;assign rom[30] = 'b001110100;assign rom[31] = 'b101010010;assign rom[32] = 'b011110111;assign rom[33] = 'b101100110;assign rom[34] = 'b010010111;assign rom[35] = 'b101100110;assign rom[36] = 'b010010111;assign rom[37] = 'b001101110;assign rom[38] = 'b001101110;assign rom[39] = 'b101000110;assign rom[40] = 'b001110100;assign rom[41] = 'b001000110;assign rom[42] = 'b001100100;assign rom[43] = 'b101100010;assign rom[44] = 'b101001100;assign rom[45] = 'b001001010;assign rom[46] = 'b111011010;assign rom[47] = 'b111011010;assign rom[48] = 'b111011010;assign rom[49] = 'b111011010;assign rom[50] = 'b111011000;assign rom[51] = 'b111011000;assign rom[52] = 'b111011000;assign rom[53] = 'b111011000;assign rom[54] = 'b101111000;assign rom[55] = 'b000110011;assign rom[56] = 'b110000010;assign rom[57] = 'b001101010;assign rom[58] = 'b001011000;assign rom[59] = 'b101001000;assign rom[60] = 'b000101011;assign rom[61] = 'b110000010;assign rom[62] = 'b111000000;assign rom[63] = 'b101001100;assign rom[64] = 'b001001010;assign rom[65] = 'b111111000;assign rom[66] = 'b111101000;assign rom[67] = 'b101001111;assign rom[68] = 'b000111010;assign rom[69] = 'b101110110;assign rom[70] = 'b101100010;assign rom[71] = 'b101001100;assign rom[72] = 'b001001010;assign rom[73] = 'b111011010;assign rom[74] = 'b111011010;assign rom[75] = 'b111011010;assign rom[76] = 'b111011010;assign rom[77] = 'b111011000;assign rom[78] = 'b111011000;assign rom[79] = 'b111011000;assign rom[80] = 'b111011000;assign rom[81] = 'b101111000;assign rom[82] = 'b000110011;assign rom[83] = 'b110000010;assign rom[84] = 'b001101010;assign rom[85] = 'b001011000;assign rom[86] = 'b101001000;assign rom[87] = 'b000101011;assign rom[88] = 'b110000010;assign rom[89] = 'b111000000;assign rom[90] = 'b101001100;assign rom[91] = 'b001001010;assign rom[92] = 'b111111000;assign rom[93] = 'b111101000;assign rom[94] = 'b101001111;assign rom[95] = 'b000111010;assign rom[96] = 'b101110110;assign rom[97] = 'b101100010;assign rom[98] = 'b101001100;assign rom[99] = 'b001001010;assign rom[100] = 'b111011010;assign rom[101] = 'b111011010;assign rom[102] = 'b111011010;assign rom[103] = 'b111011010;assign rom[104] = 'b111011000;assign rom[105] = 'b111011000;assign rom[106] = 'b111011000;assign rom[107] = 'b111011000;assign rom[108] = 'b101111000;assign rom[109] = 'b000110011;assign rom[110] = 'b110000010;assign rom[111] = 'b001101010;assign rom[112] = 'b001011000;assign rom[113] = 'b101001000;assign rom[114] = 'b000101011;assign rom[115] = 'b110000010;assign rom[116] = 'b111000000;assign rom[117] = 'b101001100;assign rom[118] = 'b001001010;assign rom[119] = 'b111111000;assign rom[120] = 'b111101000;assign rom[121] = 'b101001111;assign rom[122] = 'b000111010;assign rom[123] = 'b101110110;assign rom[124] = 'b101100010;assign rom[125] = 'b101001100;assign rom[126] = 'b001001010;assign rom[127] = 'b111011010;assign rom[128] = 'b111011010;assign rom[129] = 'b111011010;assign rom[130] = 'b111011010;assign rom[131] = 'b111011000;assign rom[132] = 'b111011000;assign rom[133] = 'b111011000;assign rom[134] = 'b111011000;assign rom[135] = 'b101111000;assign rom[136] = 'b000110011;assign rom[137] = 'b110000010;assign rom[138] = 'b001101010;assign rom[139] = 'b001011000;assign rom[140] = 'b101001000;assign rom[141] = 'b000101011;assign rom[142] = 'b110000010;assign rom[143] = 'b111000000;assign rom[144] = 'b101001100;assign rom[145] = 'b001001010;assign rom[146] = 'b111111000;assign rom[147] = 'b111101000;assign rom[148] = 'b101001111;assign rom[149] = 'b000111010;assign rom[150] = 'b101110110;assign rom[151] = 'b101100010;assign rom[152] = 'b101001100;assign rom[153] = 'b001001010;assign rom[154] = 'b111011010;assign rom[155] = 'b111011010;assign rom[156] = 'b111011010;assign rom[157] = 'b111011010;assign rom[158] = 'b111011000;assign rom[159] = 'b111011000;assign rom[160] = 'b111011000;assign rom[161] = 'b111011000;assign rom[162] = 'b101111000;assign rom[163] = 'b000110011;assign rom[164] = 'b110000010;assign rom[165] = 'b001101010;assign rom[166] = 'b001011000;assign rom[167] = 'b101001000;assign rom[168] = 'b000101011;assign rom[169] = 'b110000010;assign rom[170] = 'b111000000;assign rom[171] = 'b101001100;assign rom[172] = 'b001001010;assign rom[173] = 'b111111000;assign rom[174] = 'b111101000;assign rom[175] = 'b101001111;assign rom[176] = 'b000111010;assign rom[177] = 'b101110110;assign rom[178] = 'b101100010;assign rom[179] = 'b101001100;assign rom[180] = 'b001001010;assign rom[181] = 'b111011010;assign rom[182] = 'b111011010;assign rom[183] = 'b111011010;assign rom[184] = 'b111011010;assign rom[185] = 'b111011000;assign rom[186] = 'b111011000;assign rom[187] = 'b111011000;assign rom[188] = 'b111011000;assign rom[189] = 'b101111000;assign rom[190] = 'b000110011;assign rom[191] = 'b110000010;assign rom[192] = 'b001101010;assign rom[193] = 'b001011000;assign rom[194] = 'b101001000;assign rom[195] = 'b000101011;assign rom[196] = 'b110000010;assign rom[197] = 'b111000000;assign rom[198] = 'b101001100;assign rom[199] = 'b001001010;assign rom[200] = 'b111111000;assign rom[201] = 'b111101000;assign rom[202] = 'b101001111;assign rom[203] = 'b000111010;assign rom[204] = 'b101110110;assign rom[205] = 'b101100010;assign rom[206] = 'b101001100;assign rom[207] = 'b001001010;assign rom[208] = 'b111011010;assign rom[209] = 'b111011010;assign rom[210] = 'b111011010;assign rom[211] = 'b111011010;assign rom[212] = 'b111011000;assign rom[213] = 'b111011000;assign rom[214] = 'b111011000;assign rom[215] = 'b111011000;assign rom[216] = 'b101111000;assign rom[217] = 'b000110011;assign rom[218] = 'b110000010;assign rom[219] = 'b001101010;assign rom[220] = 'b001011000;assign rom[221] = 'b101001000;assign rom[222] = 'b000101011;assign rom[223] = 'b110000010;assign rom[224] = 'b111000000;assign rom[225] = 'b101001100;assign rom[226] = 'b001001010;assign rom[227] = 'b111111000;assign rom[228] = 'b111101000;assign rom[229] = 'b101001111;assign rom[230] = 'b000111010;assign rom[231] = 'b101110110;assign rom[232] = 'b101100010;assign rom[233] = 'b101001100;assign rom[234] = 'b001001010;assign rom[235] = 'b111011010;assign rom[236] = 'b111011010;assign rom[237] = 'b111011010;assign rom[238] = 'b111011010;assign rom[239] = 'b111011000;assign rom[240] = 'b111011000;assign rom[241] = 'b111011000;assign rom[242] = 'b111011000;assign rom[243] = 'b101111000;assign rom[244] = 'b000110011;assign rom[245] = 'b110000010;assign rom[246] = 'b001101010;assign rom[247] = 'b001011000;assign rom[248] = 'b101001000;assign rom[249] = 'b000101011;assign rom[250] = 'b110000010;assign rom[251] = 'b111000000;assign rom[252] = 'b101001100;assign rom[253] = 'b001001010;assign rom[254] = 'b111111000;assign rom[255] = 'b111101000;assign rom[256] = 'b101001111;assign rom[257] = 'b000111010;assign rom[258] = 'b101110110;assign rom[259] = 'b101100010;assign rom[260] = 'b101001100;assign rom[261] = 'b001001010;assign rom[262] = 'b111011010;assign rom[263] = 'b111011010;assign rom[264] = 'b111011010;assign rom[265] = 'b111011010;assign rom[266] = 'b111011000;assign rom[267] = 'b111011000;assign rom[268] = 'b111011000;assign rom[269] = 'b111011000;assign rom[270] = 'b101111000;assign rom[271] = 'b000110011;assign rom[272] = 'b110000010;assign rom[273] = 'b001101010;assign rom[274] = 'b001011000;assign rom[275] = 'b101001000;assign rom[276] = 'b000101011;assign rom[277] = 'b110000010;assign rom[278] = 'b111000000;assign rom[279] = 'b101001100;assign rom[280] = 'b001001010;assign rom[281] = 'b001000110;assign rom[282] = 'b001100100;assign rom[283] = 'b101100010;assign rom[284] = 'b101001100;assign rom[285] = 'b001001010;assign rom[286] = 'b111011010;assign rom[287] = 'b111011010;assign rom[288] = 'b111011010;assign rom[289] = 'b111011010;assign rom[290] = 'b111011000;assign rom[291] = 'b111011000;assign rom[292] = 'b111011000;assign rom[293] = 'b111011000;assign rom[294] = 'b101111000;assign rom[295] = 'b000110011;assign rom[296] = 'b110000010;assign rom[297] = 'b001101010;assign rom[298] = 'b001011000;assign rom[299] = 'b101001000;assign rom[300] = 'b000101011;assign rom[301] = 'b110000010;assign rom[302] = 'b111000000;assign rom[303] = 'b101001100;assign rom[304] = 'b001001010;assign rom[305] = 'b111111000;assign rom[306] = 'b111101000;assign rom[307] = 'b101001111;assign rom[308] = 'b000111010;assign rom[309] = 'b101110110;assign rom[310] = 'b101100010;assign rom[311] = 'b101001100;assign rom[312] = 'b001001010;assign rom[313] = 'b111011010;assign rom[314] = 'b111011010;assign rom[315] = 'b111011010;assign rom[316] = 'b111011010;assign rom[317] = 'b111011000;assign rom[318] = 'b111011000;assign rom[319] = 'b111011000;assign rom[320] = 'b111011000;assign rom[321] = 'b101111000;assign rom[322] = 'b000110011;assign rom[323] = 'b110000010;assign rom[324] = 'b001101010;assign rom[325] = 'b001011000;assign rom[326] = 'b101001000;assign rom[327] = 'b000101011;assign rom[328] = 'b110000010;assign rom[329] = 'b111000000;assign rom[330] = 'b101001100;assign rom[331] = 'b001001010;assign rom[332] = 'b111111000;assign rom[333] = 'b111101000;assign rom[334] = 'b101001111;assign rom[335] = 'b000111010;assign rom[336] = 'b101110110;assign rom[337] = 'b101100010;assign rom[338] = 'b101001100;assign rom[339] = 'b001001010;assign rom[340] = 'b111011010;assign rom[341] = 'b111011010;assign rom[342] = 'b111011010;assign rom[343] = 'b111011010;assign rom[344] = 'b111011000;assign rom[345] = 'b111011000;assign rom[346] = 'b111011000;assign rom[347] = 'b111011000;assign rom[348] = 'b101111000;assign rom[349] = 'b000110011;assign rom[350] = 'b110000010;assign rom[351] = 'b001101010;assign rom[352] = 'b001011000;assign rom[353] = 'b101001000;assign rom[354] = 'b000101011;assign rom[355] = 'b110000010;assign rom[356] = 'b111000000;assign rom[357] = 'b101001100;assign rom[358] = 'b001001010;assign rom[359] = 'b111111000;assign rom[360] = 'b111101000;assign rom[361] = 'b101001111;assign rom[362] = 'b000111010;assign rom[363] = 'b101110110;assign rom[364] = 'b101100010;assign rom[365] = 'b101001100;assign rom[366] = 'b001001010;assign rom[367] = 'b111011010;assign rom[368] = 'b111011010;assign rom[369] = 'b111011010;assign rom[370] = 'b111011010;assign rom[371] = 'b111011000;assign rom[372] = 'b111011000;assign rom[373] = 'b111011000;assign rom[374] = 'b111011000;assign rom[375] = 'b101111000;assign rom[376] = 'b000110011;assign rom[377] = 'b110000010;assign rom[378] = 'b001101010;assign rom[379] = 'b001011000;assign rom[380] = 'b101001000;assign rom[381] = 'b000101011;assign rom[382] = 'b110000010;assign rom[383] = 'b111000000;assign rom[384] = 'b101001100;assign rom[385] = 'b001001010;assign rom[386] = 'b111111000;assign rom[387] = 'b111101000;assign rom[388] = 'b101001111;assign rom[389] = 'b000111010;assign rom[390] = 'b101110110;assign rom[391] = 'b101100010;assign rom[392] = 'b101001100;assign rom[393] = 'b001001010;assign rom[394] = 'b111011010;assign rom[395] = 'b111011010;assign rom[396] = 'b111011010;assign rom[397] = 'b111011010;assign rom[398] = 'b111011000;assign rom[399] = 'b111011000;assign rom[400] = 'b111011000;assign rom[401] = 'b111011000;assign rom[402] = 'b101111000;assign rom[403] = 'b000110011;assign rom[404] = 'b110000010;assign rom[405] = 'b001101010;assign rom[406] = 'b001011000;assign rom[407] = 'b101001000;assign rom[408] = 'b000101011;assign rom[409] = 'b110000010;assign rom[410] = 'b111000000;assign rom[411] = 'b101001100;assign rom[412] = 'b001001010;assign rom[413] = 'b111111000;assign rom[414] = 'b111101000;assign rom[415] = 'b101001111;assign rom[416] = 'b000111010;assign rom[417] = 'b101110110;assign rom[418] = 'b101100010;assign rom[419] = 'b101001100;assign rom[420] = 'b001001010;assign rom[421] = 'b111011010;assign rom[422] = 'b111011010;assign rom[423] = 'b111011010;assign rom[424] = 'b111011010;assign rom[425] = 'b111011000;assign rom[426] = 'b111011000;assign rom[427] = 'b111011000;assign rom[428] = 'b111011000;assign rom[429] = 'b101111000;assign rom[430] = 'b000110011;assign rom[431] = 'b110000010;assign rom[432] = 'b001101010;assign rom[433] = 'b001011000;assign rom[434] = 'b101001000;assign rom[435] = 'b000101011;assign rom[436] = 'b110000010;assign rom[437] = 'b111000000;assign rom[438] = 'b101001100;assign rom[439] = 'b001001010;assign rom[440] = 'b111111000;assign rom[441] = 'b111101000;assign rom[442] = 'b101001111;assign rom[443] = 'b000111010;assign rom[444] = 'b101110110;assign rom[445] = 'b101100010;assign rom[446] = 'b101001100;assign rom[447] = 'b001001010;assign rom[448] = 'b111011010;assign rom[449] = 'b111011010;assign rom[450] = 'b111011010;assign rom[451] = 'b111011010;assign rom[452] = 'b111011000;assign rom[453] = 'b111011000;assign rom[454] = 'b111011000;assign rom[455] = 'b111011000;assign rom[456] = 'b101111000;assign rom[457] = 'b000110011;assign rom[458] = 'b110000010;assign rom[459] = 'b001101010;assign rom[460] = 'b001011000;assign rom[461] = 'b101001000;assign rom[462] = 'b000101011;assign rom[463] = 'b110000010;assign rom[464] = 'b111000000;assign rom[465] = 'b101001100;assign rom[466] = 'b001001010;assign rom[467] = 'b111111000;assign rom[468] = 'b111101000;assign rom[469] = 'b101001111;assign rom[470] = 'b000111010;assign rom[471] = 'b101110110;assign rom[472] = 'b101100010;assign rom[473] = 'b101001100;assign rom[474] = 'b001001010;assign rom[475] = 'b111011010;assign rom[476] = 'b111011010;assign rom[477] = 'b111011010;assign rom[478] = 'b111011010;assign rom[479] = 'b111011000;assign rom[480] = 'b111011000;assign rom[481] = 'b111011000;assign rom[482] = 'b111011000;assign rom[483] = 'b101111000;assign rom[484] = 'b000110011;assign rom[485] = 'b110000010;assign rom[486] = 'b001101010;assign rom[487] = 'b001011000;assign rom[488] = 'b101001000;assign rom[489] = 'b000101011;assign rom[490] = 'b110000010;assign rom[491] = 'b111000000;assign rom[492] = 'b101001100;assign rom[493] = 'b001001010;assign rom[494] = 'b111111000;assign rom[495] = 'b111101000;assign rom[496] = 'b101001111;assign rom[497] = 'b000111010;assign rom[498] = 'b101110110;assign rom[499] = 'b101100010;assign rom[500] = 'b101001100;assign rom[501] = 'b001001010;assign rom[502] = 'b111011010;assign rom[503] = 'b111011010;assign rom[504] = 'b111011010;assign rom[505] = 'b111011010;assign rom[506] = 'b111011000;assign rom[507] = 'b111011000;assign rom[508] = 'b111011000;assign rom[509] = 'b111011000;assign rom[510] = 'b101111000;assign rom[511] = 'b000110011;assign rom[512] = 'b110000010;assign rom[513] = 'b001101010;assign rom[514] = 'b001011000;assign rom[515] = 'b101001000;assign rom[516] = 'b000101011;assign rom[517] = 'b110000010;assign rom[518] = 'b111000000;assign rom[519] = 'b101001100;assign rom[520] = 'b001001010;assign rom[521] = 'b001000110;assign rom[522] = 'b001100100;assign rom[523] = 'b101100010;assign rom[524] = 'b101001100;assign rom[525] = 'b001001010;assign rom[526] = 'b111011010;assign rom[527] = 'b111011010;assign rom[528] = 'b111011010;assign rom[529] = 'b111011010;assign rom[530] = 'b111011000;assign rom[531] = 'b111011000;assign rom[532] = 'b111011000;assign rom[533] = 'b111011000;assign rom[534] = 'b101111000;assign rom[535] = 'b000110011;assign rom[536] = 'b110000010;assign rom[537] = 'b001101010;assign rom[538] = 'b001011000;assign rom[539] = 'b101001000;assign rom[540] = 'b000101011;assign rom[541] = 'b110000010;assign rom[542] = 'b111000000;assign rom[543] = 'b101001100;assign rom[544] = 'b001001010;assign rom[545] = 'b111111000;assign rom[546] = 'b111101000;assign rom[547] = 'b101001111;assign rom[548] = 'b000111010;assign rom[549] = 'b101110110;assign rom[550] = 'b101100010;assign rom[551] = 'b101001100;assign rom[552] = 'b001001010;assign rom[553] = 'b111011010;assign rom[554] = 'b111011010;assign rom[555] = 'b111011010;assign rom[556] = 'b111011010;assign rom[557] = 'b111011000;assign rom[558] = 'b111011000;assign rom[559] = 'b111011000;assign rom[560] = 'b111011000;assign rom[561] = 'b101111000;assign rom[562] = 'b000110011;assign rom[563] = 'b110000010;assign rom[564] = 'b001101010;assign rom[565] = 'b001011000;assign rom[566] = 'b101001000;assign rom[567] = 'b000101011;assign rom[568] = 'b110000010;assign rom[569] = 'b111000000;assign rom[570] = 'b101001100;assign rom[571] = 'b001001010;assign rom[572] = 'b111111000;assign rom[573] = 'b111101000;assign rom[574] = 'b101001111;assign rom[575] = 'b000111010;assign rom[576] = 'b101110110;assign rom[577] = 'b101100010;assign rom[578] = 'b101001100;assign rom[579] = 'b001001010;assign rom[580] = 'b111011010;assign rom[581] = 'b111011010;assign rom[582] = 'b111011010;assign rom[583] = 'b111011010;assign rom[584] = 'b111011000;assign rom[585] = 'b111011000;assign rom[586] = 'b111011000;assign rom[587] = 'b111011000;assign rom[588] = 'b101111000;assign rom[589] = 'b000110011;assign rom[590] = 'b110000010;assign rom[591] = 'b001101010;assign rom[592] = 'b001011000;assign rom[593] = 'b101001000;assign rom[594] = 'b000101011;assign rom[595] = 'b110000010;assign rom[596] = 'b111000000;assign rom[597] = 'b101001100;assign rom[598] = 'b001001010;assign rom[599] = 'b111111000;assign rom[600] = 'b111101000;assign rom[601] = 'b101001111;assign rom[602] = 'b000111010;assign rom[603] = 'b101110110;assign rom[604] = 'b101100010;assign rom[605] = 'b101001100;assign rom[606] = 'b001001010;assign rom[607] = 'b111011010;assign rom[608] = 'b111011010;assign rom[609] = 'b111011010;assign rom[610] = 'b111011010;assign rom[611] = 'b111011000;assign rom[612] = 'b111011000;assign rom[613] = 'b111011000;assign rom[614] = 'b111011000;assign rom[615] = 'b101111000;assign rom[616] = 'b000110011;assign rom[617] = 'b110000010;assign rom[618] = 'b001101010;assign rom[619] = 'b001011000;assign rom[620] = 'b101001000;assign rom[621] = 'b000101011;assign rom[622] = 'b110000010;assign rom[623] = 'b111000000;assign rom[624] = 'b101001100;assign rom[625] = 'b001001010;assign rom[626] = 'b111111000;assign rom[627] = 'b111101000;assign rom[628] = 'b101001111;assign rom[629] = 'b000111010;assign rom[630] = 'b101110110;assign rom[631] = 'b101100010;assign rom[632] = 'b101001100;assign rom[633] = 'b001001010;assign rom[634] = 'b111011010;assign rom[635] = 'b111011010;assign rom[636] = 'b111011010;assign rom[637] = 'b111011010;assign rom[638] = 'b111011000;assign rom[639] = 'b111011000;assign rom[640] = 'b111011000;assign rom[641] = 'b111011000;assign rom[642] = 'b101111000;assign rom[643] = 'b000110011;assign rom[644] = 'b110000010;assign rom[645] = 'b001101010;assign rom[646] = 'b001011000;assign rom[647] = 'b101001000;assign rom[648] = 'b000101011;assign rom[649] = 'b110000010;assign rom[650] = 'b111000000;assign rom[651] = 'b101001100;assign rom[652] = 'b001001010;assign rom[653] = 'b111111000;assign rom[654] = 'b111101000;assign rom[655] = 'b101001111;assign rom[656] = 'b000111010;assign rom[657] = 'b101110110;assign rom[658] = 'b101100010;assign rom[659] = 'b101001100;assign rom[660] = 'b001001010;assign rom[661] = 'b111011010;assign rom[662] = 'b111011010;assign rom[663] = 'b111011010;assign rom[664] = 'b111011010;assign rom[665] = 'b111011000;assign rom[666] = 'b111011000;assign rom[667] = 'b111011000;assign rom[668] = 'b111011000;assign rom[669] = 'b101111000;assign rom[670] = 'b000110011;assign rom[671] = 'b110000010;assign rom[672] = 'b001101010;assign rom[673] = 'b001011000;assign rom[674] = 'b101001000;assign rom[675] = 'b000101011;assign rom[676] = 'b110000010;assign rom[677] = 'b111000000;assign rom[678] = 'b101001100;assign rom[679] = 'b001001010;assign rom[680] = 'b111111000;assign rom[681] = 'b111101000;assign rom[682] = 'b101001111;assign rom[683] = 'b000111010;assign rom[684] = 'b101110110;assign rom[685] = 'b101100010;assign rom[686] = 'b101001100;assign rom[687] = 'b001001010;assign rom[688] = 'b111011010;assign rom[689] = 'b111011010;assign rom[690] = 'b111011010;assign rom[691] = 'b111011010;assign rom[692] = 'b111011000;assign rom[693] = 'b111011000;assign rom[694] = 'b111011000;assign rom[695] = 'b111011000;assign rom[696] = 'b101111000;assign rom[697] = 'b000110011;assign rom[698] = 'b110000010;assign rom[699] = 'b001101010;assign rom[700] = 'b001011000;assign rom[701] = 'b101001000;assign rom[702] = 'b000101011;assign rom[703] = 'b110000010;assign rom[704] = 'b111000000;assign rom[705] = 'b101001100;assign rom[706] = 'b001001010;assign rom[707] = 'b111111000;assign rom[708] = 'b111101000;assign rom[709] = 'b101001111;assign rom[710] = 'b000111010;assign rom[711] = 'b101110110;assign rom[712] = 'b101100010;assign rom[713] = 'b101001100;assign rom[714] = 'b001001010;assign rom[715] = 'b111011010;assign rom[716] = 'b111011010;assign rom[717] = 'b111011010;assign rom[718] = 'b111011010;assign rom[719] = 'b111011000;assign rom[720] = 'b111011000;assign rom[721] = 'b111011000;assign rom[722] = 'b111011000;assign rom[723] = 'b101111000;assign rom[724] = 'b000110011;assign rom[725] = 'b110000010;assign rom[726] = 'b001101010;assign rom[727] = 'b001011000;assign rom[728] = 'b101001000;assign rom[729] = 'b000101011;assign rom[730] = 'b110000010;assign rom[731] = 'b111000000;assign rom[732] = 'b101001100;assign rom[733] = 'b001001010;assign rom[734] = 'b111111000;assign rom[735] = 'b111101000;assign rom[736] = 'b101001111;assign rom[737] = 'b000111010;assign rom[738] = 'b101110110;assign rom[739] = 'b101100010;assign rom[740] = 'b101001100;assign rom[741] = 'b001001010;assign rom[742] = 'b111011010;assign rom[743] = 'b111011010;assign rom[744] = 'b111011010;assign rom[745] = 'b111011010;assign rom[746] = 'b111011000;assign rom[747] = 'b111011000;assign rom[748] = 'b111011000;assign rom[749] = 'b111011000;assign rom[750] = 'b101111000;assign rom[751] = 'b000110011;assign rom[752] = 'b110000010;assign rom[753] = 'b001101010;assign rom[754] = 'b001011000;assign rom[755] = 'b101001000;assign rom[756] = 'b000101011;assign rom[757] = 'b110000010;assign rom[758] = 'b111000000;assign rom[759] = 'b101001100;assign rom[760] = 'b001001010;assign rom[761] = 'b001000110;assign rom[762] = 'b001100100;assign rom[763] = 'b101100010;assign rom[764] = 'b101001100;assign rom[765] = 'b001001010;assign rom[766] = 'b111011010;assign rom[767] = 'b111011010;assign rom[768] = 'b111011010;assign rom[769] = 'b111011010;assign rom[770] = 'b111011000;assign rom[771] = 'b111011000;assign rom[772] = 'b111011000;assign rom[773] = 'b111011000;assign rom[774] = 'b101111000;assign rom[775] = 'b000110011;assign rom[776] = 'b110000010;assign rom[777] = 'b001101010;assign rom[778] = 'b001011000;assign rom[779] = 'b101001000;assign rom[780] = 'b000101011;assign rom[781] = 'b110000010;assign rom[782] = 'b111000000;assign rom[783] = 'b101001100;assign rom[784] = 'b001001010;assign rom[785] = 'b111111000;assign rom[786] = 'b111101000;assign rom[787] = 'b101001111;assign rom[788] = 'b000111010;assign rom[789] = 'b101110110;assign rom[790] = 'b101100010;assign rom[791] = 'b101001100;assign rom[792] = 'b001001010;assign rom[793] = 'b111011010;assign rom[794] = 'b111011010;assign rom[795] = 'b111011010;assign rom[796] = 'b111011010;assign rom[797] = 'b111011000;assign rom[798] = 'b111011000;assign rom[799] = 'b111011000;assign rom[800] = 'b111011000;assign rom[801] = 'b101111000;assign rom[802] = 'b000110011;assign rom[803] = 'b110000010;assign rom[804] = 'b001101010;assign rom[805] = 'b001011000;assign rom[806] = 'b101001000;assign rom[807] = 'b000101011;assign rom[808] = 'b110000010;assign rom[809] = 'b111000000;assign rom[810] = 'b101001100;assign rom[811] = 'b001001010;assign rom[812] = 'b111111000;assign rom[813] = 'b111101000;assign rom[814] = 'b101001111;assign rom[815] = 'b000111010;assign rom[816] = 'b101110110;assign rom[817] = 'b101100010;assign rom[818] = 'b101001100;assign rom[819] = 'b001001010;assign rom[820] = 'b111011010;assign rom[821] = 'b111011010;assign rom[822] = 'b111011010;assign rom[823] = 'b111011010;assign rom[824] = 'b111011000;assign rom[825] = 'b111011000;assign rom[826] = 'b111011000;assign rom[827] = 'b111011000;assign rom[828] = 'b101111000;assign rom[829] = 'b000110011;assign rom[830] = 'b110000010;assign rom[831] = 'b001101010;assign rom[832] = 'b001011000;assign rom[833] = 'b101001000;assign rom[834] = 'b000101011;assign rom[835] = 'b110000010;assign rom[836] = 'b111000000;assign rom[837] = 'b101001100;assign rom[838] = 'b001001010;assign rom[839] = 'b111111000;assign rom[840] = 'b111101000;assign rom[841] = 'b101001111;assign rom[842] = 'b000111010;assign rom[843] = 'b101110110;assign rom[844] = 'b101100010;assign rom[845] = 'b101001100;assign rom[846] = 'b001001010;assign rom[847] = 'b111011010;assign rom[848] = 'b111011010;assign rom[849] = 'b111011010;assign rom[850] = 'b111011010;assign rom[851] = 'b111011000;assign rom[852] = 'b111011000;assign rom[853] = 'b111011000;assign rom[854] = 'b111011000;assign rom[855] = 'b101111000;assign rom[856] = 'b000110011;assign rom[857] = 'b110000010;assign rom[858] = 'b001101010;assign rom[859] = 'b001011000;assign rom[860] = 'b101001000;assign rom[861] = 'b000101011;assign rom[862] = 'b110000010;assign rom[863] = 'b111000000;assign rom[864] = 'b101001100;assign rom[865] = 'b001001010;assign rom[866] = 'b111111000;assign rom[867] = 'b111101000;assign rom[868] = 'b101001111;assign rom[869] = 'b000111010;assign rom[870] = 'b101110110;assign rom[871] = 'b101100010;assign rom[872] = 'b101001100;assign rom[873] = 'b001001010;assign rom[874] = 'b111011010;assign rom[875] = 'b111011010;assign rom[876] = 'b111011010;assign rom[877] = 'b111011010;assign rom[878] = 'b111011000;assign rom[879] = 'b111011000;assign rom[880] = 'b111011000;assign rom[881] = 'b111011000;assign rom[882] = 'b101111000;assign rom[883] = 'b000110011;assign rom[884] = 'b110000010;assign rom[885] = 'b001101010;assign rom[886] = 'b001011000;assign rom[887] = 'b101001000;assign rom[888] = 'b000101011;assign rom[889] = 'b110000010;assign rom[890] = 'b111000000;assign rom[891] = 'b101001100;assign rom[892] = 'b001001010;assign rom[893] = 'b111111000;assign rom[894] = 'b111101000;assign rom[895] = 'b101001111;assign rom[896] = 'b000111010;assign rom[897] = 'b101110110;assign rom[898] = 'b101100010;assign rom[899] = 'b101001100;assign rom[900] = 'b001001010;assign rom[901] = 'b111011010;assign rom[902] = 'b111011010;assign rom[903] = 'b111011010;assign rom[904] = 'b111011010;assign rom[905] = 'b111011000;assign rom[906] = 'b111011000;assign rom[907] = 'b111011000;assign rom[908] = 'b111011000;assign rom[909] = 'b101111000;assign rom[910] = 'b000110011;assign rom[911] = 'b110000010;assign rom[912] = 'b001101010;assign rom[913] = 'b001011000;assign rom[914] = 'b101001000;assign rom[915] = 'b000101011;assign rom[916] = 'b110000010;assign rom[917] = 'b111000000;assign rom[918] = 'b101001100;assign rom[919] = 'b001001010;assign rom[920] = 'b111111000;assign rom[921] = 'b111101000;assign rom[922] = 'b101001111;assign rom[923] = 'b000111010;assign rom[924] = 'b101110110;assign rom[925] = 'b101100010;assign rom[926] = 'b101001100;assign rom[927] = 'b001001010;assign rom[928] = 'b111011010;assign rom[929] = 'b111011010;assign rom[930] = 'b111011010;assign rom[931] = 'b111011010;assign rom[932] = 'b111011000;assign rom[933] = 'b111011000;assign rom[934] = 'b111011000;assign rom[935] = 'b111011000;assign rom[936] = 'b101111000;assign rom[937] = 'b000110011;assign rom[938] = 'b110000010;assign rom[939] = 'b001101010;assign rom[940] = 'b001011000;assign rom[941] = 'b101001000;assign rom[942] = 'b000101011;assign rom[943] = 'b110000010;assign rom[944] = 'b111000000;assign rom[945] = 'b101001100;assign rom[946] = 'b001001010;assign rom[947] = 'b111111000;assign rom[948] = 'b111101000;assign rom[949] = 'b101001111;assign rom[950] = 'b000111010;assign rom[951] = 'b101110110;assign rom[952] = 'b101100010;assign rom[953] = 'b101001100;assign rom[954] = 'b001001010;assign rom[955] = 'b111011010;assign rom[956] = 'b111011010;assign rom[957] = 'b111011010;assign rom[958] = 'b111011010;assign rom[959] = 'b111011000;assign rom[960] = 'b111011000;assign rom[961] = 'b111011000;assign rom[962] = 'b111011000;assign rom[963] = 'b101111000;assign rom[964] = 'b000110011;assign rom[965] = 'b110000010;assign rom[966] = 'b001101010;assign rom[967] = 'b001011000;assign rom[968] = 'b101001000;assign rom[969] = 'b000101011;assign rom[970] = 'b110000010;assign rom[971] = 'b111000000;assign rom[972] = 'b101001100;assign rom[973] = 'b001001010;assign rom[974] = 'b111111000;assign rom[975] = 'b111101000;assign rom[976] = 'b101001111;assign rom[977] = 'b000111010;assign rom[978] = 'b101110110;assign rom[979] = 'b101100010;assign rom[980] = 'b101001100;assign rom[981] = 'b001001010;assign rom[982] = 'b111011010;assign rom[983] = 'b111011010;assign rom[984] = 'b111011010;assign rom[985] = 'b111011010;assign rom[986] = 'b111011000;assign rom[987] = 'b111011000;assign rom[988] = 'b111011000;assign rom[989] = 'b111011000;assign rom[990] = 'b101111000;assign rom[991] = 'b000110011;assign rom[992] = 'b110000010;assign rom[993] = 'b001101010;assign rom[994] = 'b001011000;assign rom[995] = 'b101001000;assign rom[996] = 'b000101011;assign rom[997] = 'b110000010;assign rom[998] = 'b111000000;assign rom[999] = 'b101001100;assign rom[1000] = 'b001001010;assign rom[1001] = 'b001000110;assign rom[1002] = 'b001100100;assign rom[1003] = 'b101100010;assign rom[1004] = 'b101001100;assign rom[1005] = 'b001001010;assign rom[1006] = 'b111011010;assign rom[1007] = 'b111011010;assign rom[1008] = 'b111011010;assign rom[1009] = 'b111011010;assign rom[1010] = 'b111011000;assign rom[1011] = 'b111011000;assign rom[1012] = 'b111011000;assign rom[1013] = 'b111011000;assign rom[1014] = 'b101111000;assign rom[1015] = 'b000110011;assign rom[1016] = 'b110000010;assign rom[1017] = 'b001101010;assign rom[1018] = 'b001011000;assign rom[1019] = 'b101001000;assign rom[1020] = 'b000101011;assign rom[1021] = 'b110000010;assign rom[1022] = 'b111000000;assign rom[1023] = 'b101001100;assign rom[1024] = 'b001001010;assign rom[1025] = 'b111111000;assign rom[1026] = 'b111101000;assign rom[1027] = 'b101001111;assign rom[1028] = 'b000111010;assign rom[1029] = 'b101110110;assign rom[1030] = 'b101100010;assign rom[1031] = 'b101001100;assign rom[1032] = 'b001001010;assign rom[1033] = 'b111011010;assign rom[1034] = 'b111011010;assign rom[1035] = 'b111011010;assign rom[1036] = 'b111011010;assign rom[1037] = 'b111011000;assign rom[1038] = 'b111011000;assign rom[1039] = 'b111011000;assign rom[1040] = 'b111011000;assign rom[1041] = 'b101111000;assign rom[1042] = 'b000110011;assign rom[1043] = 'b110000010;assign rom[1044] = 'b001101010;assign rom[1045] = 'b001011000;assign rom[1046] = 'b101001000;assign rom[1047] = 'b000101011;assign rom[1048] = 'b110000010;assign rom[1049] = 'b111000000;assign rom[1050] = 'b101001100;assign rom[1051] = 'b001001010;assign rom[1052] = 'b111111000;assign rom[1053] = 'b111101000;assign rom[1054] = 'b101001111;assign rom[1055] = 'b000111010;assign rom[1056] = 'b101110110;assign rom[1057] = 'b101100010;assign rom[1058] = 'b101001100;assign rom[1059] = 'b001001010;assign rom[1060] = 'b111011010;assign rom[1061] = 'b111011010;assign rom[1062] = 'b111011010;assign rom[1063] = 'b111011010;assign rom[1064] = 'b111011000;assign rom[1065] = 'b111011000;assign rom[1066] = 'b111011000;assign rom[1067] = 'b111011000;assign rom[1068] = 'b101111000;assign rom[1069] = 'b000110011;assign rom[1070] = 'b110000010;assign rom[1071] = 'b001101010;assign rom[1072] = 'b001011000;assign rom[1073] = 'b101001000;assign rom[1074] = 'b000101011;assign rom[1075] = 'b110000010;assign rom[1076] = 'b111000000;assign rom[1077] = 'b101001100;assign rom[1078] = 'b001001010;assign rom[1079] = 'b111111000;assign rom[1080] = 'b111101000;assign rom[1081] = 'b101001111;assign rom[1082] = 'b000111010;assign rom[1083] = 'b101110110;assign rom[1084] = 'b101100010;assign rom[1085] = 'b101001100;assign rom[1086] = 'b001001010;assign rom[1087] = 'b111011010;assign rom[1088] = 'b111011010;assign rom[1089] = 'b111011010;assign rom[1090] = 'b111011010;assign rom[1091] = 'b111011000;assign rom[1092] = 'b111011000;assign rom[1093] = 'b111011000;assign rom[1094] = 'b111011000;assign rom[1095] = 'b101111000;assign rom[1096] = 'b000110011;assign rom[1097] = 'b110000010;assign rom[1098] = 'b001101010;assign rom[1099] = 'b001011000;assign rom[1100] = 'b101001000;assign rom[1101] = 'b000101011;assign rom[1102] = 'b110000010;assign rom[1103] = 'b111000000;assign rom[1104] = 'b101001100;assign rom[1105] = 'b001001010;assign rom[1106] = 'b111111000;assign rom[1107] = 'b111101000;assign rom[1108] = 'b101001111;assign rom[1109] = 'b000111010;assign rom[1110] = 'b101110110;assign rom[1111] = 'b101100010;assign rom[1112] = 'b101001100;assign rom[1113] = 'b001001010;assign rom[1114] = 'b111011010;assign rom[1115] = 'b111011010;assign rom[1116] = 'b111011010;assign rom[1117] = 'b111011010;assign rom[1118] = 'b111011000;assign rom[1119] = 'b111011000;assign rom[1120] = 'b111011000;assign rom[1121] = 'b111011000;assign rom[1122] = 'b101111000;assign rom[1123] = 'b000110011;assign rom[1124] = 'b110000010;assign rom[1125] = 'b001101010;assign rom[1126] = 'b001011000;assign rom[1127] = 'b101001000;assign rom[1128] = 'b000101011;assign rom[1129] = 'b110000010;assign rom[1130] = 'b111000000;assign rom[1131] = 'b101001100;assign rom[1132] = 'b001001010;assign rom[1133] = 'b111111000;assign rom[1134] = 'b111101000;assign rom[1135] = 'b101001111;assign rom[1136] = 'b000111010;assign rom[1137] = 'b101110110;assign rom[1138] = 'b101100010;assign rom[1139] = 'b101001100;assign rom[1140] = 'b001001010;assign rom[1141] = 'b111011010;assign rom[1142] = 'b111011010;assign rom[1143] = 'b111011010;assign rom[1144] = 'b111011010;assign rom[1145] = 'b111011000;assign rom[1146] = 'b111011000;assign rom[1147] = 'b111011000;assign rom[1148] = 'b111011000;assign rom[1149] = 'b101111000;assign rom[1150] = 'b000110011;assign rom[1151] = 'b110000010;assign rom[1152] = 'b001101010;assign rom[1153] = 'b001011000;assign rom[1154] = 'b101001000;assign rom[1155] = 'b000101011;assign rom[1156] = 'b110000010;assign rom[1157] = 'b111000000;assign rom[1158] = 'b101001100;assign rom[1159] = 'b001001010;assign rom[1160] = 'b111111000;assign rom[1161] = 'b111101000;assign rom[1162] = 'b101001111;assign rom[1163] = 'b000111010;assign rom[1164] = 'b101110110;assign rom[1165] = 'b101100010;assign rom[1166] = 'b101001100;assign rom[1167] = 'b001001010;assign rom[1168] = 'b111011010;assign rom[1169] = 'b111011010;assign rom[1170] = 'b111011010;assign rom[1171] = 'b111011010;assign rom[1172] = 'b111011000;assign rom[1173] = 'b111011000;assign rom[1174] = 'b111011000;assign rom[1175] = 'b111011000;assign rom[1176] = 'b101111000;assign rom[1177] = 'b000110011;assign rom[1178] = 'b110000010;assign rom[1179] = 'b001101010;assign rom[1180] = 'b001011000;assign rom[1181] = 'b101001000;assign rom[1182] = 'b000101011;assign rom[1183] = 'b110000010;assign rom[1184] = 'b111000000;assign rom[1185] = 'b101001100;assign rom[1186] = 'b001001010;assign rom[1187] = 'b111111000;assign rom[1188] = 'b111101000;assign rom[1189] = 'b101001111;assign rom[1190] = 'b000111010;assign rom[1191] = 'b101110110;assign rom[1192] = 'b101100010;assign rom[1193] = 'b101001100;assign rom[1194] = 'b001001010;assign rom[1195] = 'b111011010;assign rom[1196] = 'b111011010;assign rom[1197] = 'b111011010;assign rom[1198] = 'b111011010;assign rom[1199] = 'b111011000;assign rom[1200] = 'b111011000;assign rom[1201] = 'b111011000;assign rom[1202] = 'b111011000;assign rom[1203] = 'b101111000;assign rom[1204] = 'b000110011;assign rom[1205] = 'b110000010;assign rom[1206] = 'b001101010;assign rom[1207] = 'b001011000;assign rom[1208] = 'b101001000;assign rom[1209] = 'b000101011;assign rom[1210] = 'b110000010;assign rom[1211] = 'b111000000;assign rom[1212] = 'b101001100;assign rom[1213] = 'b001001010;assign rom[1214] = 'b111111000;assign rom[1215] = 'b111101000;assign rom[1216] = 'b101001111;assign rom[1217] = 'b000111010;assign rom[1218] = 'b101110110;assign rom[1219] = 'b101100010;assign rom[1220] = 'b101001100;assign rom[1221] = 'b001001010;assign rom[1222] = 'b111011010;assign rom[1223] = 'b111011010;assign rom[1224] = 'b111011010;assign rom[1225] = 'b111011010;assign rom[1226] = 'b111011000;assign rom[1227] = 'b111011000;assign rom[1228] = 'b111011000;assign rom[1229] = 'b111011000;assign rom[1230] = 'b101111000;assign rom[1231] = 'b000110011;assign rom[1232] = 'b110000010;assign rom[1233] = 'b001101010;assign rom[1234] = 'b001011000;assign rom[1235] = 'b101001000;assign rom[1236] = 'b000101011;assign rom[1237] = 'b110000010;assign rom[1238] = 'b111000000;assign rom[1239] = 'b101001100;assign rom[1240] = 'b001001010;assign rom[1241] = 'b001000110;assign rom[1242] = 'b001100100;assign rom[1243] = 'b101100010;assign rom[1244] = 'b101001100;assign rom[1245] = 'b001001010;assign rom[1246] = 'b111011010;assign rom[1247] = 'b111011010;assign rom[1248] = 'b111011010;assign rom[1249] = 'b111011010;assign rom[1250] = 'b111011000;assign rom[1251] = 'b111011000;assign rom[1252] = 'b111011000;assign rom[1253] = 'b111011000;assign rom[1254] = 'b101111000;assign rom[1255] = 'b000110011;assign rom[1256] = 'b110000010;assign rom[1257] = 'b001101010;assign rom[1258] = 'b001011000;assign rom[1259] = 'b101001000;assign rom[1260] = 'b000101011;assign rom[1261] = 'b110000010;assign rom[1262] = 'b111000000;assign rom[1263] = 'b101001100;assign rom[1264] = 'b001001010;assign rom[1265] = 'b111111000;assign rom[1266] = 'b111101000;assign rom[1267] = 'b101001111;assign rom[1268] = 'b000111010;assign rom[1269] = 'b101110110;assign rom[1270] = 'b101100010;assign rom[1271] = 'b101001100;assign rom[1272] = 'b001001010;assign rom[1273] = 'b111011010;assign rom[1274] = 'b111011010;assign rom[1275] = 'b111011010;assign rom[1276] = 'b111011010;assign rom[1277] = 'b111011000;assign rom[1278] = 'b111011000;assign rom[1279] = 'b111011000;assign rom[1280] = 'b111011000;assign rom[1281] = 'b101111000;assign rom[1282] = 'b000110011;assign rom[1283] = 'b110000010;assign rom[1284] = 'b001101010;assign rom[1285] = 'b001011000;assign rom[1286] = 'b101001000;assign rom[1287] = 'b000101011;assign rom[1288] = 'b110000010;assign rom[1289] = 'b111000000;assign rom[1290] = 'b101001100;assign rom[1291] = 'b001001010;assign rom[1292] = 'b111111000;assign rom[1293] = 'b111101000;assign rom[1294] = 'b101001111;assign rom[1295] = 'b000111010;assign rom[1296] = 'b101110110;assign rom[1297] = 'b101100010;assign rom[1298] = 'b101001100;assign rom[1299] = 'b001001010;assign rom[1300] = 'b111011010;assign rom[1301] = 'b111011010;assign rom[1302] = 'b111011010;assign rom[1303] = 'b111011010;assign rom[1304] = 'b111011000;assign rom[1305] = 'b111011000;assign rom[1306] = 'b111011000;assign rom[1307] = 'b111011000;assign rom[1308] = 'b101111000;assign rom[1309] = 'b000110011;assign rom[1310] = 'b110000010;assign rom[1311] = 'b001101010;assign rom[1312] = 'b001011000;assign rom[1313] = 'b101001000;assign rom[1314] = 'b000101011;assign rom[1315] = 'b110000010;assign rom[1316] = 'b111000000;assign rom[1317] = 'b101001100;assign rom[1318] = 'b001001010;assign rom[1319] = 'b111111000;assign rom[1320] = 'b111101000;assign rom[1321] = 'b101001111;assign rom[1322] = 'b000111010;assign rom[1323] = 'b101110110;assign rom[1324] = 'b101100010;assign rom[1325] = 'b101001100;assign rom[1326] = 'b001001010;assign rom[1327] = 'b111011010;assign rom[1328] = 'b111011010;assign rom[1329] = 'b111011010;assign rom[1330] = 'b111011010;assign rom[1331] = 'b111011000;assign rom[1332] = 'b111011000;assign rom[1333] = 'b111011000;assign rom[1334] = 'b111011000;assign rom[1335] = 'b101111000;assign rom[1336] = 'b000110011;assign rom[1337] = 'b110000010;assign rom[1338] = 'b001101010;assign rom[1339] = 'b001011000;assign rom[1340] = 'b101001000;assign rom[1341] = 'b000101011;assign rom[1342] = 'b110000010;assign rom[1343] = 'b111000000;assign rom[1344] = 'b101001100;assign rom[1345] = 'b001001010;assign rom[1346] = 'b111111000;assign rom[1347] = 'b111101000;assign rom[1348] = 'b101001111;assign rom[1349] = 'b000111010;assign rom[1350] = 'b101110110;assign rom[1351] = 'b101100010;assign rom[1352] = 'b101001100;assign rom[1353] = 'b001001010;assign rom[1354] = 'b111011010;assign rom[1355] = 'b111011010;assign rom[1356] = 'b111011010;assign rom[1357] = 'b111011010;assign rom[1358] = 'b111011000;assign rom[1359] = 'b111011000;assign rom[1360] = 'b111011000;assign rom[1361] = 'b111011000;assign rom[1362] = 'b101111000;assign rom[1363] = 'b000110011;assign rom[1364] = 'b110000010;assign rom[1365] = 'b001101010;assign rom[1366] = 'b001011000;assign rom[1367] = 'b101001000;assign rom[1368] = 'b000101011;assign rom[1369] = 'b110000010;assign rom[1370] = 'b111000000;assign rom[1371] = 'b101001100;assign rom[1372] = 'b001001010;assign rom[1373] = 'b111111000;assign rom[1374] = 'b111101000;assign rom[1375] = 'b101001111;assign rom[1376] = 'b000111010;assign rom[1377] = 'b101110110;assign rom[1378] = 'b101100010;assign rom[1379] = 'b101001100;assign rom[1380] = 'b001001010;assign rom[1381] = 'b111011010;assign rom[1382] = 'b111011010;assign rom[1383] = 'b111011010;assign rom[1384] = 'b111011010;assign rom[1385] = 'b111011000;assign rom[1386] = 'b111011000;assign rom[1387] = 'b111011000;assign rom[1388] = 'b111011000;assign rom[1389] = 'b101111000;assign rom[1390] = 'b000110011;assign rom[1391] = 'b110000010;assign rom[1392] = 'b001101010;assign rom[1393] = 'b001011000;assign rom[1394] = 'b101001000;assign rom[1395] = 'b000101011;assign rom[1396] = 'b110000010;assign rom[1397] = 'b111000000;assign rom[1398] = 'b101001100;assign rom[1399] = 'b001001010;assign rom[1400] = 'b111111000;assign rom[1401] = 'b111101000;assign rom[1402] = 'b101001111;assign rom[1403] = 'b000111010;assign rom[1404] = 'b101110110;assign rom[1405] = 'b101100010;assign rom[1406] = 'b101001100;assign rom[1407] = 'b001001010;assign rom[1408] = 'b111011010;assign rom[1409] = 'b111011010;assign rom[1410] = 'b111011010;assign rom[1411] = 'b111011010;assign rom[1412] = 'b111011000;assign rom[1413] = 'b111011000;assign rom[1414] = 'b111011000;assign rom[1415] = 'b111011000;assign rom[1416] = 'b101111000;assign rom[1417] = 'b000110011;assign rom[1418] = 'b110000010;assign rom[1419] = 'b001101010;assign rom[1420] = 'b001011000;assign rom[1421] = 'b101001000;assign rom[1422] = 'b000101011;assign rom[1423] = 'b110000010;assign rom[1424] = 'b111000000;assign rom[1425] = 'b101001100;assign rom[1426] = 'b001001010;assign rom[1427] = 'b111111000;assign rom[1428] = 'b111101000;assign rom[1429] = 'b101001111;assign rom[1430] = 'b000111010;assign rom[1431] = 'b101110110;assign rom[1432] = 'b101100010;assign rom[1433] = 'b101001100;assign rom[1434] = 'b001001010;assign rom[1435] = 'b111011010;assign rom[1436] = 'b111011010;assign rom[1437] = 'b111011010;assign rom[1438] = 'b111011010;assign rom[1439] = 'b111011000;assign rom[1440] = 'b111011000;assign rom[1441] = 'b111011000;assign rom[1442] = 'b111011000;assign rom[1443] = 'b101111000;assign rom[1444] = 'b000110011;assign rom[1445] = 'b110000010;assign rom[1446] = 'b001101010;assign rom[1447] = 'b001011000;assign rom[1448] = 'b101001000;assign rom[1449] = 'b000101011;assign rom[1450] = 'b110000010;assign rom[1451] = 'b111000000;assign rom[1452] = 'b101001100;assign rom[1453] = 'b001001010;assign rom[1454] = 'b111111000;assign rom[1455] = 'b111101000;assign rom[1456] = 'b101001111;assign rom[1457] = 'b000111010;assign rom[1458] = 'b101110110;assign rom[1459] = 'b101100010;assign rom[1460] = 'b101001100;assign rom[1461] = 'b001001010;assign rom[1462] = 'b111011010;assign rom[1463] = 'b111011010;assign rom[1464] = 'b111011010;assign rom[1465] = 'b111011010;assign rom[1466] = 'b111011000;assign rom[1467] = 'b111011000;assign rom[1468] = 'b111011000;assign rom[1469] = 'b111011000;assign rom[1470] = 'b101111000;assign rom[1471] = 'b000110011;assign rom[1472] = 'b110000010;assign rom[1473] = 'b001101010;assign rom[1474] = 'b001011000;assign rom[1475] = 'b101001000;assign rom[1476] = 'b000101011;assign rom[1477] = 'b110000010;assign rom[1478] = 'b111000000;assign rom[1479] = 'b101001100;assign rom[1480] = 'b001001010;assign rom[1481] = 'b001000110;assign rom[1482] = 'b001100100;assign rom[1483] = 'b101100010;assign rom[1484] = 'b101001100;assign rom[1485] = 'b001001010;assign rom[1486] = 'b111011010;assign rom[1487] = 'b111011010;assign rom[1488] = 'b111011010;assign rom[1489] = 'b111011010;assign rom[1490] = 'b111011000;assign rom[1491] = 'b111011000;assign rom[1492] = 'b111011000;assign rom[1493] = 'b111011000;assign rom[1494] = 'b101111000;assign rom[1495] = 'b000110011;assign rom[1496] = 'b110000010;assign rom[1497] = 'b001101010;assign rom[1498] = 'b001011000;assign rom[1499] = 'b101001000;assign rom[1500] = 'b000101011;assign rom[1501] = 'b110000010;assign rom[1502] = 'b111000000;assign rom[1503] = 'b101001100;assign rom[1504] = 'b001001010;assign rom[1505] = 'b111111000;assign rom[1506] = 'b111101000;assign rom[1507] = 'b101001111;assign rom[1508] = 'b000111010;assign rom[1509] = 'b101110110;assign rom[1510] = 'b101100010;assign rom[1511] = 'b101001100;assign rom[1512] = 'b001001010;assign rom[1513] = 'b111011010;assign rom[1514] = 'b111011010;assign rom[1515] = 'b111011010;assign rom[1516] = 'b111011010;assign rom[1517] = 'b111011000;assign rom[1518] = 'b111011000;assign rom[1519] = 'b111011000;assign rom[1520] = 'b111011000;assign rom[1521] = 'b101111000;assign rom[1522] = 'b000110011;assign rom[1523] = 'b110000010;assign rom[1524] = 'b001101010;assign rom[1525] = 'b001011000;assign rom[1526] = 'b101001000;assign rom[1527] = 'b000101011;assign rom[1528] = 'b110000010;assign rom[1529] = 'b111000000;assign rom[1530] = 'b101001100;assign rom[1531] = 'b001001010;assign rom[1532] = 'b111111000;assign rom[1533] = 'b111101000;assign rom[1534] = 'b101001111;assign rom[1535] = 'b000111010;assign rom[1536] = 'b101110110;assign rom[1537] = 'b101100010;assign rom[1538] = 'b101001100;assign rom[1539] = 'b001001010;assign rom[1540] = 'b111011010;assign rom[1541] = 'b111011010;assign rom[1542] = 'b111011010;assign rom[1543] = 'b111011010;assign rom[1544] = 'b111011000;assign rom[1545] = 'b111011000;assign rom[1546] = 'b111011000;assign rom[1547] = 'b111011000;assign rom[1548] = 'b101111000;assign rom[1549] = 'b000110011;assign rom[1550] = 'b110000010;assign rom[1551] = 'b001101010;assign rom[1552] = 'b001011000;assign rom[1553] = 'b101001000;assign rom[1554] = 'b000101011;assign rom[1555] = 'b110000010;assign rom[1556] = 'b111000000;assign rom[1557] = 'b101001100;assign rom[1558] = 'b001001010;assign rom[1559] = 'b111111000;assign rom[1560] = 'b111101000;assign rom[1561] = 'b101001111;assign rom[1562] = 'b000111010;assign rom[1563] = 'b101110110;assign rom[1564] = 'b101100010;assign rom[1565] = 'b101001100;assign rom[1566] = 'b001001010;assign rom[1567] = 'b111011010;assign rom[1568] = 'b111011010;assign rom[1569] = 'b111011010;assign rom[1570] = 'b111011010;assign rom[1571] = 'b111011000;assign rom[1572] = 'b111011000;assign rom[1573] = 'b111011000;assign rom[1574] = 'b111011000;assign rom[1575] = 'b101111000;assign rom[1576] = 'b000110011;assign rom[1577] = 'b110000010;assign rom[1578] = 'b001101010;assign rom[1579] = 'b001011000;assign rom[1580] = 'b101001000;assign rom[1581] = 'b000101011;assign rom[1582] = 'b110000010;assign rom[1583] = 'b111000000;assign rom[1584] = 'b101001100;assign rom[1585] = 'b001001010;assign rom[1586] = 'b111111000;assign rom[1587] = 'b111101000;assign rom[1588] = 'b101001111;assign rom[1589] = 'b000111010;assign rom[1590] = 'b101110110;assign rom[1591] = 'b101100010;assign rom[1592] = 'b101001100;assign rom[1593] = 'b001001010;assign rom[1594] = 'b111011010;assign rom[1595] = 'b111011010;assign rom[1596] = 'b111011010;assign rom[1597] = 'b111011010;assign rom[1598] = 'b111011000;assign rom[1599] = 'b111011000;assign rom[1600] = 'b111011000;assign rom[1601] = 'b111011000;assign rom[1602] = 'b101111000;assign rom[1603] = 'b000110011;assign rom[1604] = 'b110000010;assign rom[1605] = 'b001101010;assign rom[1606] = 'b001011000;assign rom[1607] = 'b101001000;assign rom[1608] = 'b000101011;assign rom[1609] = 'b110000010;assign rom[1610] = 'b111000000;assign rom[1611] = 'b101001100;assign rom[1612] = 'b001001010;assign rom[1613] = 'b111111000;assign rom[1614] = 'b111101000;assign rom[1615] = 'b101001111;assign rom[1616] = 'b000111010;assign rom[1617] = 'b101110110;assign rom[1618] = 'b101100010;assign rom[1619] = 'b101001100;assign rom[1620] = 'b001001010;assign rom[1621] = 'b111011010;assign rom[1622] = 'b111011010;assign rom[1623] = 'b111011010;assign rom[1624] = 'b111011010;assign rom[1625] = 'b111011000;assign rom[1626] = 'b111011000;assign rom[1627] = 'b111011000;assign rom[1628] = 'b111011000;assign rom[1629] = 'b101111000;assign rom[1630] = 'b000110011;assign rom[1631] = 'b110000010;assign rom[1632] = 'b001101010;assign rom[1633] = 'b001011000;assign rom[1634] = 'b101001000;assign rom[1635] = 'b000101011;assign rom[1636] = 'b110000010;assign rom[1637] = 'b111000000;assign rom[1638] = 'b101001100;assign rom[1639] = 'b001001010;assign rom[1640] = 'b111111000;assign rom[1641] = 'b111101000;assign rom[1642] = 'b101001111;assign rom[1643] = 'b000111010;assign rom[1644] = 'b101110110;assign rom[1645] = 'b101100010;assign rom[1646] = 'b101001100;assign rom[1647] = 'b001001010;assign rom[1648] = 'b111011010;assign rom[1649] = 'b111011010;assign rom[1650] = 'b111011010;assign rom[1651] = 'b111011010;assign rom[1652] = 'b111011000;assign rom[1653] = 'b111011000;assign rom[1654] = 'b111011000;assign rom[1655] = 'b111011000;assign rom[1656] = 'b101111000;assign rom[1657] = 'b000110011;assign rom[1658] = 'b110000010;assign rom[1659] = 'b001101010;assign rom[1660] = 'b001011000;assign rom[1661] = 'b101001000;assign rom[1662] = 'b000101011;assign rom[1663] = 'b110000010;assign rom[1664] = 'b111000000;assign rom[1665] = 'b101001100;assign rom[1666] = 'b001001010;assign rom[1667] = 'b111111000;assign rom[1668] = 'b111101000;assign rom[1669] = 'b101001111;assign rom[1670] = 'b000111010;assign rom[1671] = 'b101110110;assign rom[1672] = 'b101100010;assign rom[1673] = 'b101001100;assign rom[1674] = 'b001001010;assign rom[1675] = 'b111011010;assign rom[1676] = 'b111011010;assign rom[1677] = 'b111011010;assign rom[1678] = 'b111011010;assign rom[1679] = 'b111011000;assign rom[1680] = 'b111011000;assign rom[1681] = 'b111011000;assign rom[1682] = 'b111011000;assign rom[1683] = 'b101111000;assign rom[1684] = 'b000110011;assign rom[1685] = 'b110000010;assign rom[1686] = 'b001101010;assign rom[1687] = 'b001011000;assign rom[1688] = 'b101001000;assign rom[1689] = 'b000101011;assign rom[1690] = 'b110000010;assign rom[1691] = 'b111000000;assign rom[1692] = 'b101001100;assign rom[1693] = 'b001001010;assign rom[1694] = 'b111111000;assign rom[1695] = 'b111101000;assign rom[1696] = 'b101001111;assign rom[1697] = 'b000111010;assign rom[1698] = 'b101110110;assign rom[1699] = 'b101100010;assign rom[1700] = 'b101001100;assign rom[1701] = 'b001001010;assign rom[1702] = 'b111011010;assign rom[1703] = 'b111011010;assign rom[1704] = 'b111011010;assign rom[1705] = 'b111011010;assign rom[1706] = 'b111011000;assign rom[1707] = 'b111011000;assign rom[1708] = 'b111011000;assign rom[1709] = 'b111011000;assign rom[1710] = 'b101111000;assign rom[1711] = 'b000110011;assign rom[1712] = 'b110000010;assign rom[1713] = 'b001101010;assign rom[1714] = 'b001011000;assign rom[1715] = 'b101001000;assign rom[1716] = 'b000101011;assign rom[1717] = 'b110000010;assign rom[1718] = 'b111000000;assign rom[1719] = 'b101001100;assign rom[1720] = 'b001001010;assign rom[1721] = 'b001000110;assign rom[1722] = 'b001100100;assign rom[1723] = 'b101100010;assign rom[1724] = 'b101001100;assign rom[1725] = 'b001001010;assign rom[1726] = 'b111011010;assign rom[1727] = 'b111011010;assign rom[1728] = 'b111011010;assign rom[1729] = 'b111011010;assign rom[1730] = 'b111011000;assign rom[1731] = 'b111011000;assign rom[1732] = 'b111011000;assign rom[1733] = 'b111011000;assign rom[1734] = 'b101111000;assign rom[1735] = 'b000110011;assign rom[1736] = 'b110000010;assign rom[1737] = 'b001101010;assign rom[1738] = 'b001011000;assign rom[1739] = 'b101001000;assign rom[1740] = 'b000101011;assign rom[1741] = 'b110000010;assign rom[1742] = 'b111000000;assign rom[1743] = 'b101001100;assign rom[1744] = 'b001001010;assign rom[1745] = 'b111111000;assign rom[1746] = 'b111101000;assign rom[1747] = 'b101001111;assign rom[1748] = 'b000111010;assign rom[1749] = 'b101110110;assign rom[1750] = 'b101100010;assign rom[1751] = 'b101001100;assign rom[1752] = 'b001001010;assign rom[1753] = 'b111011010;assign rom[1754] = 'b111011010;assign rom[1755] = 'b111011010;assign rom[1756] = 'b111011010;assign rom[1757] = 'b111011000;assign rom[1758] = 'b111011000;assign rom[1759] = 'b111011000;assign rom[1760] = 'b111011000;assign rom[1761] = 'b101111000;assign rom[1762] = 'b000110011;assign rom[1763] = 'b110000010;assign rom[1764] = 'b001101010;assign rom[1765] = 'b001011000;assign rom[1766] = 'b101001000;assign rom[1767] = 'b000101011;assign rom[1768] = 'b110000010;assign rom[1769] = 'b111000000;assign rom[1770] = 'b101001100;assign rom[1771] = 'b001001010;assign rom[1772] = 'b111111000;assign rom[1773] = 'b111101000;assign rom[1774] = 'b101001111;assign rom[1775] = 'b000111010;assign rom[1776] = 'b101110110;assign rom[1777] = 'b101100010;assign rom[1778] = 'b101001100;assign rom[1779] = 'b001001010;assign rom[1780] = 'b111011010;assign rom[1781] = 'b111011010;assign rom[1782] = 'b111011010;assign rom[1783] = 'b111011010;assign rom[1784] = 'b111011000;assign rom[1785] = 'b111011000;assign rom[1786] = 'b111011000;assign rom[1787] = 'b111011000;assign rom[1788] = 'b101111000;assign rom[1789] = 'b000110011;assign rom[1790] = 'b110000010;assign rom[1791] = 'b001101010;assign rom[1792] = 'b001011000;assign rom[1793] = 'b101001000;assign rom[1794] = 'b000101011;assign rom[1795] = 'b110000010;assign rom[1796] = 'b111000000;assign rom[1797] = 'b101001100;assign rom[1798] = 'b001001010;assign rom[1799] = 'b111111000;assign rom[1800] = 'b111101000;assign rom[1801] = 'b101001111;assign rom[1802] = 'b000111010;assign rom[1803] = 'b101110110;assign rom[1804] = 'b101100010;assign rom[1805] = 'b101001100;assign rom[1806] = 'b001001010;assign rom[1807] = 'b111011010;assign rom[1808] = 'b111011010;assign rom[1809] = 'b111011010;assign rom[1810] = 'b111011010;assign rom[1811] = 'b111011000;assign rom[1812] = 'b111011000;assign rom[1813] = 'b111011000;assign rom[1814] = 'b111011000;assign rom[1815] = 'b101111000;assign rom[1816] = 'b000110011;assign rom[1817] = 'b110000010;assign rom[1818] = 'b001101010;assign rom[1819] = 'b001011000;assign rom[1820] = 'b101001000;assign rom[1821] = 'b000101011;assign rom[1822] = 'b110000010;assign rom[1823] = 'b111000000;assign rom[1824] = 'b101001100;assign rom[1825] = 'b001001010;assign rom[1826] = 'b111111000;assign rom[1827] = 'b111101000;assign rom[1828] = 'b101001111;assign rom[1829] = 'b000111010;assign rom[1830] = 'b101110110;assign rom[1831] = 'b101100010;assign rom[1832] = 'b101001100;assign rom[1833] = 'b001001010;assign rom[1834] = 'b111011010;assign rom[1835] = 'b111011010;assign rom[1836] = 'b111011010;assign rom[1837] = 'b111011010;assign rom[1838] = 'b111011000;assign rom[1839] = 'b111011000;assign rom[1840] = 'b111011000;assign rom[1841] = 'b111011000;assign rom[1842] = 'b101111000;assign rom[1843] = 'b000110011;assign rom[1844] = 'b110000010;assign rom[1845] = 'b001101010;assign rom[1846] = 'b001011000;assign rom[1847] = 'b101001000;assign rom[1848] = 'b000101011;assign rom[1849] = 'b110000010;assign rom[1850] = 'b111000000;assign rom[1851] = 'b101001100;assign rom[1852] = 'b001001010;assign rom[1853] = 'b111111000;assign rom[1854] = 'b111101000;assign rom[1855] = 'b101001111;assign rom[1856] = 'b000111010;assign rom[1857] = 'b101110110;assign rom[1858] = 'b101100010;assign rom[1859] = 'b101001100;assign rom[1860] = 'b001001010;assign rom[1861] = 'b111011010;assign rom[1862] = 'b111011010;assign rom[1863] = 'b111011010;assign rom[1864] = 'b111011010;assign rom[1865] = 'b111011000;assign rom[1866] = 'b111011000;assign rom[1867] = 'b111011000;assign rom[1868] = 'b111011000;assign rom[1869] = 'b101111000;assign rom[1870] = 'b000110011;assign rom[1871] = 'b110000010;assign rom[1872] = 'b001101010;assign rom[1873] = 'b001011000;assign rom[1874] = 'b101001000;assign rom[1875] = 'b000101011;assign rom[1876] = 'b110000010;assign rom[1877] = 'b111000000;assign rom[1878] = 'b101001100;assign rom[1879] = 'b001001010;assign rom[1880] = 'b111111000;assign rom[1881] = 'b111101000;assign rom[1882] = 'b101001111;assign rom[1883] = 'b000111010;assign rom[1884] = 'b101110110;assign rom[1885] = 'b101100010;assign rom[1886] = 'b101001100;assign rom[1887] = 'b001001010;assign rom[1888] = 'b111011010;assign rom[1889] = 'b111011010;assign rom[1890] = 'b111011010;assign rom[1891] = 'b111011010;assign rom[1892] = 'b111011000;assign rom[1893] = 'b111011000;assign rom[1894] = 'b111011000;assign rom[1895] = 'b111011000;assign rom[1896] = 'b101111000;assign rom[1897] = 'b000110011;assign rom[1898] = 'b110000010;assign rom[1899] = 'b001101010;assign rom[1900] = 'b001011000;assign rom[1901] = 'b101001000;assign rom[1902] = 'b000101011;assign rom[1903] = 'b110000010;assign rom[1904] = 'b111000000;assign rom[1905] = 'b101001100;assign rom[1906] = 'b001001010;assign rom[1907] = 'b111111000;assign rom[1908] = 'b111101000;assign rom[1909] = 'b101001111;assign rom[1910] = 'b000111010;assign rom[1911] = 'b101110110;assign rom[1912] = 'b101100010;assign rom[1913] = 'b101001100;assign rom[1914] = 'b001001010;assign rom[1915] = 'b111011010;assign rom[1916] = 'b111011010;assign rom[1917] = 'b111011010;assign rom[1918] = 'b111011010;assign rom[1919] = 'b111011000;assign rom[1920] = 'b111011000;assign rom[1921] = 'b111011000;assign rom[1922] = 'b111011000;assign rom[1923] = 'b101111000;assign rom[1924] = 'b000110011;assign rom[1925] = 'b110000010;assign rom[1926] = 'b001101010;assign rom[1927] = 'b001011000;assign rom[1928] = 'b101001000;assign rom[1929] = 'b000101011;assign rom[1930] = 'b110000010;assign rom[1931] = 'b111000000;assign rom[1932] = 'b101001100;assign rom[1933] = 'b001001010;assign rom[1934] = 'b111111000;assign rom[1935] = 'b111101000;assign rom[1936] = 'b101001111;assign rom[1937] = 'b000111010;assign rom[1938] = 'b101110110;assign rom[1939] = 'b101100010;assign rom[1940] = 'b101001100;assign rom[1941] = 'b001001010;assign rom[1942] = 'b111011010;assign rom[1943] = 'b111011010;assign rom[1944] = 'b111011010;assign rom[1945] = 'b111011010;assign rom[1946] = 'b111011000;assign rom[1947] = 'b111011000;assign rom[1948] = 'b111011000;assign rom[1949] = 'b111011000;assign rom[1950] = 'b101111000;assign rom[1951] = 'b000110011;assign rom[1952] = 'b110000010;assign rom[1953] = 'b001101010;assign rom[1954] = 'b001011000;assign rom[1955] = 'b101001000;assign rom[1956] = 'b000101011;assign rom[1957] = 'b110000010;assign rom[1958] = 'b111000000;assign rom[1959] = 'b101001100;assign rom[1960] = 'b001001010;assign rom[1961] = 'b001000110;assign rom[1962] = 'b001100100;assign rom[1963] = 'b101100010;assign rom[1964] = 'b101001100;assign rom[1965] = 'b001001010;assign rom[1966] = 'b111011010;assign rom[1967] = 'b111011010;assign rom[1968] = 'b111011010;assign rom[1969] = 'b111011010;assign rom[1970] = 'b111011000;assign rom[1971] = 'b111011000;assign rom[1972] = 'b111011000;assign rom[1973] = 'b111011000;assign rom[1974] = 'b101111000;assign rom[1975] = 'b000110011;assign rom[1976] = 'b110000010;assign rom[1977] = 'b001101010;assign rom[1978] = 'b001011000;assign rom[1979] = 'b101001000;assign rom[1980] = 'b000101011;assign rom[1981] = 'b110000010;assign rom[1982] = 'b111000000;assign rom[1983] = 'b101001100;assign rom[1984] = 'b001001010;assign rom[1985] = 'b111111000;assign rom[1986] = 'b111101000;assign rom[1987] = 'b101001111;assign rom[1988] = 'b000111010;assign rom[1989] = 'b101110110;assign rom[1990] = 'b101100010;assign rom[1991] = 'b101001100;assign rom[1992] = 'b001001010;assign rom[1993] = 'b111011010;assign rom[1994] = 'b111011010;assign rom[1995] = 'b111011010;assign rom[1996] = 'b111011010;assign rom[1997] = 'b111011000;assign rom[1998] = 'b111011000;assign rom[1999] = 'b111011000;assign rom[2000] = 'b111011000;assign rom[2001] = 'b101111000;assign rom[2002] = 'b000110011;assign rom[2003] = 'b110000010;assign rom[2004] = 'b001101010;assign rom[2005] = 'b001011000;assign rom[2006] = 'b101001000;assign rom[2007] = 'b000101011;assign rom[2008] = 'b110000010;assign rom[2009] = 'b111000000;assign rom[2010] = 'b101001100;assign rom[2011] = 'b001001010;assign rom[2012] = 'b111111000;assign rom[2013] = 'b111101000;assign rom[2014] = 'b101001111;assign rom[2015] = 'b000111010;assign rom[2016] = 'b101110110;assign rom[2017] = 'b101100010;assign rom[2018] = 'b101001100;assign rom[2019] = 'b001001010;assign rom[2020] = 'b111011010;assign rom[2021] = 'b111011010;assign rom[2022] = 'b111011010;assign rom[2023] = 'b111011010;assign rom[2024] = 'b111011000;assign rom[2025] = 'b111011000;assign rom[2026] = 'b111011000;assign rom[2027] = 'b111011000;assign rom[2028] = 'b101111000;assign rom[2029] = 'b000110011;assign rom[2030] = 'b110000010;assign rom[2031] = 'b001101010;assign rom[2032] = 'b001011000;assign rom[2033] = 'b101001000;assign rom[2034] = 'b000101011;assign rom[2035] = 'b110000010;assign rom[2036] = 'b111000000;assign rom[2037] = 'b101001100;assign rom[2038] = 'b001001010;assign rom[2039] = 'b111111000;assign rom[2040] = 'b111101000;assign rom[2041] = 'b101001111;assign rom[2042] = 'b000111010;assign rom[2043] = 'b101110110;assign rom[2044] = 'b101100010;assign rom[2045] = 'b101001100;assign rom[2046] = 'b001001010;assign rom[2047] = 'b111011010;assign rom[2048] = 'b111011010;assign rom[2049] = 'b111011010;assign rom[2050] = 'b111011010;assign rom[2051] = 'b111011000;assign rom[2052] = 'b111011000;assign rom[2053] = 'b111011000;assign rom[2054] = 'b111011000;assign rom[2055] = 'b101111000;assign rom[2056] = 'b000110011;assign rom[2057] = 'b110000010;assign rom[2058] = 'b001101010;assign rom[2059] = 'b001011000;assign rom[2060] = 'b101001000;assign rom[2061] = 'b000101011;assign rom[2062] = 'b110000010;assign rom[2063] = 'b111000000;assign rom[2064] = 'b101001100;assign rom[2065] = 'b001001010;assign rom[2066] = 'b111111000;assign rom[2067] = 'b111101000;assign rom[2068] = 'b101001111;assign rom[2069] = 'b000111010;assign rom[2070] = 'b101110110;assign rom[2071] = 'b101100010;assign rom[2072] = 'b101001100;assign rom[2073] = 'b001001010;assign rom[2074] = 'b111011010;assign rom[2075] = 'b111011010;assign rom[2076] = 'b111011010;assign rom[2077] = 'b111011010;assign rom[2078] = 'b111011000;assign rom[2079] = 'b111011000;assign rom[2080] = 'b111011000;assign rom[2081] = 'b111011000;assign rom[2082] = 'b101111000;assign rom[2083] = 'b000110011;assign rom[2084] = 'b110000010;assign rom[2085] = 'b001101010;assign rom[2086] = 'b001011000;assign rom[2087] = 'b101001000;assign rom[2088] = 'b000101011;assign rom[2089] = 'b110000010;assign rom[2090] = 'b111000000;assign rom[2091] = 'b101001100;assign rom[2092] = 'b001001010;assign rom[2093] = 'b111111000;assign rom[2094] = 'b111101000;assign rom[2095] = 'b101001111;assign rom[2096] = 'b000111010;assign rom[2097] = 'b101110110;assign rom[2098] = 'b101100010;assign rom[2099] = 'b101001100;assign rom[2100] = 'b001001010;assign rom[2101] = 'b111011010;assign rom[2102] = 'b111011010;assign rom[2103] = 'b111011010;assign rom[2104] = 'b111011010;assign rom[2105] = 'b111011000;assign rom[2106] = 'b111011000;assign rom[2107] = 'b111011000;assign rom[2108] = 'b111011000;assign rom[2109] = 'b101111000;assign rom[2110] = 'b000110011;assign rom[2111] = 'b110000010;assign rom[2112] = 'b001101010;assign rom[2113] = 'b001011000;assign rom[2114] = 'b101001000;assign rom[2115] = 'b000101011;assign rom[2116] = 'b110000010;assign rom[2117] = 'b111000000;assign rom[2118] = 'b101001100;assign rom[2119] = 'b001001010;assign rom[2120] = 'b111111000;assign rom[2121] = 'b111101000;assign rom[2122] = 'b101001111;assign rom[2123] = 'b000111010;assign rom[2124] = 'b101110110;assign rom[2125] = 'b101100010;assign rom[2126] = 'b101001100;assign rom[2127] = 'b001001010;assign rom[2128] = 'b111011010;assign rom[2129] = 'b111011010;assign rom[2130] = 'b111011010;assign rom[2131] = 'b111011010;assign rom[2132] = 'b111011000;assign rom[2133] = 'b111011000;assign rom[2134] = 'b111011000;assign rom[2135] = 'b111011000;assign rom[2136] = 'b101111000;assign rom[2137] = 'b000110011;assign rom[2138] = 'b110000010;assign rom[2139] = 'b001101010;assign rom[2140] = 'b001011000;assign rom[2141] = 'b101001000;assign rom[2142] = 'b000101011;assign rom[2143] = 'b110000010;assign rom[2144] = 'b111000000;assign rom[2145] = 'b101001100;assign rom[2146] = 'b001001010;assign rom[2147] = 'b111111000;assign rom[2148] = 'b111101000;assign rom[2149] = 'b101001111;assign rom[2150] = 'b000111010;assign rom[2151] = 'b101110110;assign rom[2152] = 'b101100010;assign rom[2153] = 'b101001100;assign rom[2154] = 'b001001010;assign rom[2155] = 'b111011010;assign rom[2156] = 'b111011010;assign rom[2157] = 'b111011010;assign rom[2158] = 'b111011010;assign rom[2159] = 'b111011000;assign rom[2160] = 'b111011000;assign rom[2161] = 'b111011000;assign rom[2162] = 'b111011000;assign rom[2163] = 'b101111000;assign rom[2164] = 'b000110011;assign rom[2165] = 'b110000010;assign rom[2166] = 'b001101010;assign rom[2167] = 'b001011000;assign rom[2168] = 'b101001000;assign rom[2169] = 'b000101011;assign rom[2170] = 'b110000010;assign rom[2171] = 'b111000000;assign rom[2172] = 'b101001100;assign rom[2173] = 'b001001010;assign rom[2174] = 'b111111000;assign rom[2175] = 'b111101000;assign rom[2176] = 'b101001111;assign rom[2177] = 'b000111010;assign rom[2178] = 'b101110110;assign rom[2179] = 'b101100010;assign rom[2180] = 'b101001100;assign rom[2181] = 'b001001010;assign rom[2182] = 'b111011010;assign rom[2183] = 'b111011010;assign rom[2184] = 'b111011010;assign rom[2185] = 'b111011010;assign rom[2186] = 'b111011000;assign rom[2187] = 'b111011000;assign rom[2188] = 'b111011000;assign rom[2189] = 'b111011000;assign rom[2190] = 'b101111000;assign rom[2191] = 'b000110011;assign rom[2192] = 'b110000010;assign rom[2193] = 'b001101010;assign rom[2194] = 'b001011000;assign rom[2195] = 'b101001000;assign rom[2196] = 'b000101011;assign rom[2197] = 'b110000010;assign rom[2198] = 'b111000000;assign rom[2199] = 'b101001100;assign rom[2200] = 'b001001010;assign rom[2201] = 'b001000110;assign rom[2202] = 'b001100100;assign rom[2203] = 'b101100010;assign rom[2204] = 'b101001100;assign rom[2205] = 'b001001010;assign rom[2206] = 'b111011010;assign rom[2207] = 'b111011010;assign rom[2208] = 'b111011010;assign rom[2209] = 'b111011010;assign rom[2210] = 'b111011000;assign rom[2211] = 'b111011000;assign rom[2212] = 'b111011000;assign rom[2213] = 'b111011000;assign rom[2214] = 'b101111000;assign rom[2215] = 'b000110011;assign rom[2216] = 'b110000010;assign rom[2217] = 'b001101010;assign rom[2218] = 'b001011000;assign rom[2219] = 'b101001000;assign rom[2220] = 'b000101011;assign rom[2221] = 'b110000010;assign rom[2222] = 'b111000000;assign rom[2223] = 'b101001100;assign rom[2224] = 'b001001010;assign rom[2225] = 'b111111000;assign rom[2226] = 'b111101000;assign rom[2227] = 'b101001111;assign rom[2228] = 'b000111010;assign rom[2229] = 'b101110110;assign rom[2230] = 'b101100010;assign rom[2231] = 'b101001100;assign rom[2232] = 'b001001010;assign rom[2233] = 'b111011010;assign rom[2234] = 'b111011010;assign rom[2235] = 'b111011010;assign rom[2236] = 'b111011010;assign rom[2237] = 'b111011000;assign rom[2238] = 'b111011000;assign rom[2239] = 'b111011000;assign rom[2240] = 'b111011000;assign rom[2241] = 'b101111000;assign rom[2242] = 'b000110011;assign rom[2243] = 'b110000010;assign rom[2244] = 'b001101010;assign rom[2245] = 'b001011000;assign rom[2246] = 'b101001000;assign rom[2247] = 'b000101011;assign rom[2248] = 'b110000010;assign rom[2249] = 'b111000000;assign rom[2250] = 'b101001100;assign rom[2251] = 'b001001010;assign rom[2252] = 'b111111000;assign rom[2253] = 'b111101000;assign rom[2254] = 'b101001111;assign rom[2255] = 'b000111010;assign rom[2256] = 'b101110110;assign rom[2257] = 'b101100010;assign rom[2258] = 'b101001100;assign rom[2259] = 'b001001010;assign rom[2260] = 'b111011010;assign rom[2261] = 'b111011010;assign rom[2262] = 'b111011010;assign rom[2263] = 'b111011010;assign rom[2264] = 'b111011000;assign rom[2265] = 'b111011000;assign rom[2266] = 'b111011000;assign rom[2267] = 'b111011000;assign rom[2268] = 'b101111000;assign rom[2269] = 'b000110011;assign rom[2270] = 'b110000010;assign rom[2271] = 'b001101010;assign rom[2272] = 'b001011000;assign rom[2273] = 'b101001000;assign rom[2274] = 'b000101011;assign rom[2275] = 'b110000010;assign rom[2276] = 'b111000000;assign rom[2277] = 'b101001100;assign rom[2278] = 'b001001010;assign rom[2279] = 'b111111000;assign rom[2280] = 'b111101000;assign rom[2281] = 'b101001111;assign rom[2282] = 'b000111010;assign rom[2283] = 'b101110110;assign rom[2284] = 'b101100010;assign rom[2285] = 'b101001100;assign rom[2286] = 'b001001010;assign rom[2287] = 'b111011010;assign rom[2288] = 'b111011010;assign rom[2289] = 'b111011010;assign rom[2290] = 'b111011010;assign rom[2291] = 'b111011000;assign rom[2292] = 'b111011000;assign rom[2293] = 'b111011000;assign rom[2294] = 'b111011000;assign rom[2295] = 'b101111000;assign rom[2296] = 'b000110011;assign rom[2297] = 'b110000010;assign rom[2298] = 'b001101010;assign rom[2299] = 'b001011000;assign rom[2300] = 'b101001000;assign rom[2301] = 'b000101011;assign rom[2302] = 'b110000010;assign rom[2303] = 'b111000000;assign rom[2304] = 'b101001100;assign rom[2305] = 'b001001010;assign rom[2306] = 'b111111000;assign rom[2307] = 'b111101000;assign rom[2308] = 'b101001111;assign rom[2309] = 'b000111010;assign rom[2310] = 'b101110110;assign rom[2311] = 'b101100010;assign rom[2312] = 'b101001100;assign rom[2313] = 'b001001010;assign rom[2314] = 'b111011010;assign rom[2315] = 'b111011010;assign rom[2316] = 'b111011010;assign rom[2317] = 'b111011010;assign rom[2318] = 'b111011000;assign rom[2319] = 'b111011000;assign rom[2320] = 'b111011000;assign rom[2321] = 'b111011000;assign rom[2322] = 'b101111000;assign rom[2323] = 'b000110011;assign rom[2324] = 'b110000010;assign rom[2325] = 'b001101010;assign rom[2326] = 'b001011000;assign rom[2327] = 'b101001000;assign rom[2328] = 'b000101011;assign rom[2329] = 'b110000010;assign rom[2330] = 'b111000000;assign rom[2331] = 'b101001100;assign rom[2332] = 'b001001010;assign rom[2333] = 'b111111000;assign rom[2334] = 'b111101000;assign rom[2335] = 'b101001111;assign rom[2336] = 'b000111010;assign rom[2337] = 'b101110110;assign rom[2338] = 'b101100010;assign rom[2339] = 'b101001100;assign rom[2340] = 'b001001010;assign rom[2341] = 'b111011010;assign rom[2342] = 'b111011010;assign rom[2343] = 'b111011010;assign rom[2344] = 'b111011010;assign rom[2345] = 'b111011000;assign rom[2346] = 'b111011000;assign rom[2347] = 'b111011000;assign rom[2348] = 'b111011000;assign rom[2349] = 'b101111000;assign rom[2350] = 'b000110011;assign rom[2351] = 'b110000010;assign rom[2352] = 'b001101010;assign rom[2353] = 'b001011000;assign rom[2354] = 'b101001000;assign rom[2355] = 'b000101011;assign rom[2356] = 'b110000010;assign rom[2357] = 'b111000000;assign rom[2358] = 'b101001100;assign rom[2359] = 'b001001010;assign rom[2360] = 'b111111000;assign rom[2361] = 'b111101000;assign rom[2362] = 'b101001111;assign rom[2363] = 'b000111010;assign rom[2364] = 'b101110110;assign rom[2365] = 'b101100010;assign rom[2366] = 'b101001100;assign rom[2367] = 'b001001010;assign rom[2368] = 'b111011010;assign rom[2369] = 'b111011010;assign rom[2370] = 'b111011010;assign rom[2371] = 'b111011010;assign rom[2372] = 'b111011000;assign rom[2373] = 'b111011000;assign rom[2374] = 'b111011000;assign rom[2375] = 'b111011000;assign rom[2376] = 'b101111000;assign rom[2377] = 'b000110011;assign rom[2378] = 'b110000010;assign rom[2379] = 'b001101010;assign rom[2380] = 'b001011000;assign rom[2381] = 'b101001000;assign rom[2382] = 'b000101011;assign rom[2383] = 'b110000010;assign rom[2384] = 'b111000000;assign rom[2385] = 'b101001100;assign rom[2386] = 'b001001010;assign rom[2387] = 'b111111000;assign rom[2388] = 'b111101000;assign rom[2389] = 'b101001111;assign rom[2390] = 'b000111010;assign rom[2391] = 'b101110110;assign rom[2392] = 'b101100010;assign rom[2393] = 'b101001100;assign rom[2394] = 'b001001010;assign rom[2395] = 'b111011010;assign rom[2396] = 'b111011010;assign rom[2397] = 'b111011010;assign rom[2398] = 'b111011010;assign rom[2399] = 'b111011000;assign rom[2400] = 'b111011000;assign rom[2401] = 'b111011000;assign rom[2402] = 'b111011000;assign rom[2403] = 'b101111000;assign rom[2404] = 'b000110011;assign rom[2405] = 'b110000010;assign rom[2406] = 'b001101010;assign rom[2407] = 'b001011000;assign rom[2408] = 'b101001000;assign rom[2409] = 'b000101011;assign rom[2410] = 'b110000010;assign rom[2411] = 'b111000000;assign rom[2412] = 'b101001100;assign rom[2413] = 'b001001010;assign rom[2414] = 'b111111000;assign rom[2415] = 'b111101000;assign rom[2416] = 'b101001111;assign rom[2417] = 'b000111010;assign rom[2418] = 'b101110110;assign rom[2419] = 'b101100010;assign rom[2420] = 'b101001100;assign rom[2421] = 'b001001010;assign rom[2422] = 'b111011010;assign rom[2423] = 'b111011010;assign rom[2424] = 'b111011010;assign rom[2425] = 'b111011010;assign rom[2426] = 'b111011000;assign rom[2427] = 'b111011000;assign rom[2428] = 'b111011000;assign rom[2429] = 'b111011000;assign rom[2430] = 'b101111000;assign rom[2431] = 'b000110011;assign rom[2432] = 'b110000010;assign rom[2433] = 'b001101010;assign rom[2434] = 'b001011000;assign rom[2435] = 'b101001000;assign rom[2436] = 'b000101011;assign rom[2437] = 'b110000010;assign rom[2438] = 'b111000000;assign rom[2439] = 'b101001100;assign rom[2440] = 'b001001010;assign rom[2441] = 'b001000110;assign rom[2442] = 'b001100100;assign rom[2443] = 'b101100010;assign rom[2444] = 'b101001100;assign rom[2445] = 'b001001010;assign rom[2446] = 'b111011010;assign rom[2447] = 'b111011010;assign rom[2448] = 'b111011010;assign rom[2449] = 'b111011010;assign rom[2450] = 'b111011000;assign rom[2451] = 'b111011000;assign rom[2452] = 'b111011000;assign rom[2453] = 'b111011000;assign rom[2454] = 'b101111000;assign rom[2455] = 'b000110011;assign rom[2456] = 'b110000010;assign rom[2457] = 'b001101010;assign rom[2458] = 'b001011000;assign rom[2459] = 'b101001000;assign rom[2460] = 'b000101011;assign rom[2461] = 'b110000010;assign rom[2462] = 'b111000000;assign rom[2463] = 'b101001100;assign rom[2464] = 'b001001010;assign rom[2465] = 'b111111000;assign rom[2466] = 'b111101000;assign rom[2467] = 'b101001111;assign rom[2468] = 'b000111010;assign rom[2469] = 'b101110110;assign rom[2470] = 'b101100010;assign rom[2471] = 'b101001100;assign rom[2472] = 'b001001010;assign rom[2473] = 'b111011010;assign rom[2474] = 'b111011010;assign rom[2475] = 'b111011010;assign rom[2476] = 'b111011010;assign rom[2477] = 'b111011000;assign rom[2478] = 'b111011000;assign rom[2479] = 'b111011000;assign rom[2480] = 'b111011000;assign rom[2481] = 'b101111000;assign rom[2482] = 'b000110011;assign rom[2483] = 'b110000010;assign rom[2484] = 'b001101010;assign rom[2485] = 'b001011000;assign rom[2486] = 'b101001000;assign rom[2487] = 'b000101011;assign rom[2488] = 'b110000010;assign rom[2489] = 'b111000000;assign rom[2490] = 'b101001100;assign rom[2491] = 'b001001010;assign rom[2492] = 'b111111000;assign rom[2493] = 'b111101000;assign rom[2494] = 'b101001111;assign rom[2495] = 'b000111010;assign rom[2496] = 'b101110110;assign rom[2497] = 'b101100010;assign rom[2498] = 'b101001100;assign rom[2499] = 'b001001010;assign rom[2500] = 'b111011010;assign rom[2501] = 'b111011010;assign rom[2502] = 'b111011010;assign rom[2503] = 'b111011010;assign rom[2504] = 'b111011000;assign rom[2505] = 'b111011000;assign rom[2506] = 'b111011000;assign rom[2507] = 'b111011000;assign rom[2508] = 'b101111000;assign rom[2509] = 'b000110011;assign rom[2510] = 'b110000010;assign rom[2511] = 'b001101010;assign rom[2512] = 'b001011000;assign rom[2513] = 'b101001000;assign rom[2514] = 'b000101011;assign rom[2515] = 'b110000010;assign rom[2516] = 'b111000000;assign rom[2517] = 'b101001100;assign rom[2518] = 'b001001010;assign rom[2519] = 'b111111000;assign rom[2520] = 'b111101000;assign rom[2521] = 'b101001111;assign rom[2522] = 'b000111010;assign rom[2523] = 'b101110110;assign rom[2524] = 'b101100010;assign rom[2525] = 'b101001100;assign rom[2526] = 'b001001010;assign rom[2527] = 'b111011010;assign rom[2528] = 'b111011010;assign rom[2529] = 'b111011010;assign rom[2530] = 'b111011010;assign rom[2531] = 'b111011000;assign rom[2532] = 'b111011000;assign rom[2533] = 'b111011000;assign rom[2534] = 'b111011000;assign rom[2535] = 'b101111000;assign rom[2536] = 'b000110011;assign rom[2537] = 'b110000010;assign rom[2538] = 'b001101010;assign rom[2539] = 'b001011000;assign rom[2540] = 'b101001000;assign rom[2541] = 'b000101011;assign rom[2542] = 'b110000010;assign rom[2543] = 'b111000000;assign rom[2544] = 'b101001100;assign rom[2545] = 'b001001010;assign rom[2546] = 'b111111000;assign rom[2547] = 'b111101000;assign rom[2548] = 'b101001111;assign rom[2549] = 'b000111010;assign rom[2550] = 'b101110110;assign rom[2551] = 'b101100010;assign rom[2552] = 'b101001100;assign rom[2553] = 'b001001010;assign rom[2554] = 'b111011010;assign rom[2555] = 'b111011010;assign rom[2556] = 'b111011010;assign rom[2557] = 'b111011010;assign rom[2558] = 'b111011000;assign rom[2559] = 'b111011000;assign rom[2560] = 'b111011000;assign rom[2561] = 'b111011000;assign rom[2562] = 'b101111000;assign rom[2563] = 'b000110011;assign rom[2564] = 'b110000010;assign rom[2565] = 'b001101010;assign rom[2566] = 'b001011000;assign rom[2567] = 'b101001000;assign rom[2568] = 'b000101011;assign rom[2569] = 'b110000010;assign rom[2570] = 'b111000000;assign rom[2571] = 'b101001100;assign rom[2572] = 'b001001010;assign rom[2573] = 'b111111000;assign rom[2574] = 'b111101000;assign rom[2575] = 'b101001111;assign rom[2576] = 'b000111010;assign rom[2577] = 'b101110110;assign rom[2578] = 'b101100010;assign rom[2579] = 'b101001100;assign rom[2580] = 'b001001010;assign rom[2581] = 'b111011010;assign rom[2582] = 'b111011010;assign rom[2583] = 'b111011010;assign rom[2584] = 'b111011010;assign rom[2585] = 'b111011000;assign rom[2586] = 'b111011000;assign rom[2587] = 'b111011000;assign rom[2588] = 'b111011000;assign rom[2589] = 'b101111000;assign rom[2590] = 'b000110011;assign rom[2591] = 'b110000010;assign rom[2592] = 'b001101010;assign rom[2593] = 'b001011000;assign rom[2594] = 'b101001000;assign rom[2595] = 'b000101011;assign rom[2596] = 'b110000010;assign rom[2597] = 'b111000000;assign rom[2598] = 'b101001100;assign rom[2599] = 'b001001010;assign rom[2600] = 'b111111000;assign rom[2601] = 'b111101000;assign rom[2602] = 'b101001111;assign rom[2603] = 'b000111010;assign rom[2604] = 'b101110110;assign rom[2605] = 'b101100010;assign rom[2606] = 'b101001100;assign rom[2607] = 'b001001010;assign rom[2608] = 'b111011010;assign rom[2609] = 'b111011010;assign rom[2610] = 'b111011010;assign rom[2611] = 'b111011010;assign rom[2612] = 'b111011000;assign rom[2613] = 'b111011000;assign rom[2614] = 'b111011000;assign rom[2615] = 'b111011000;assign rom[2616] = 'b101111000;assign rom[2617] = 'b000110011;assign rom[2618] = 'b110000010;assign rom[2619] = 'b001101010;assign rom[2620] = 'b001011000;assign rom[2621] = 'b101001000;assign rom[2622] = 'b000101011;assign rom[2623] = 'b110000010;assign rom[2624] = 'b111000000;assign rom[2625] = 'b101001100;assign rom[2626] = 'b001001010;assign rom[2627] = 'b111111000;assign rom[2628] = 'b111101000;assign rom[2629] = 'b101001111;assign rom[2630] = 'b000111010;assign rom[2631] = 'b101110110;assign rom[2632] = 'b101100010;assign rom[2633] = 'b101001100;assign rom[2634] = 'b001001010;assign rom[2635] = 'b111011010;assign rom[2636] = 'b111011010;assign rom[2637] = 'b111011010;assign rom[2638] = 'b111011010;assign rom[2639] = 'b111011000;assign rom[2640] = 'b111011000;assign rom[2641] = 'b111011000;assign rom[2642] = 'b111011000;assign rom[2643] = 'b101111000;assign rom[2644] = 'b000110011;assign rom[2645] = 'b110000010;assign rom[2646] = 'b001101010;assign rom[2647] = 'b001011000;assign rom[2648] = 'b101001000;assign rom[2649] = 'b000101011;assign rom[2650] = 'b110000010;assign rom[2651] = 'b111000000;assign rom[2652] = 'b101001100;assign rom[2653] = 'b001001010;assign rom[2654] = 'b111111000;assign rom[2655] = 'b111101000;assign rom[2656] = 'b101001111;assign rom[2657] = 'b000111010;assign rom[2658] = 'b101110110;assign rom[2659] = 'b101100010;assign rom[2660] = 'b101001100;assign rom[2661] = 'b001001010;assign rom[2662] = 'b111011010;assign rom[2663] = 'b111011010;assign rom[2664] = 'b111011010;assign rom[2665] = 'b111011010;assign rom[2666] = 'b111011000;assign rom[2667] = 'b111011000;assign rom[2668] = 'b111011000;assign rom[2669] = 'b111011000;assign rom[2670] = 'b101111000;assign rom[2671] = 'b000110011;assign rom[2672] = 'b110000010;assign rom[2673] = 'b001101010;assign rom[2674] = 'b001011000;assign rom[2675] = 'b101001000;assign rom[2676] = 'b000101011;assign rom[2677] = 'b110000010;assign rom[2678] = 'b111000000;assign rom[2679] = 'b101001100;assign rom[2680] = 'b001001010;assign rom[2681] = 'b001000110;assign rom[2682] = 'b001100100;assign rom[2683] = 'b101100010;assign rom[2684] = 'b101001100;assign rom[2685] = 'b001001010;assign rom[2686] = 'b111011010;assign rom[2687] = 'b111011010;assign rom[2688] = 'b111011010;assign rom[2689] = 'b111011010;assign rom[2690] = 'b111011000;assign rom[2691] = 'b111011000;assign rom[2692] = 'b111011000;assign rom[2693] = 'b111011000;assign rom[2694] = 'b101111000;assign rom[2695] = 'b000110011;assign rom[2696] = 'b110000010;assign rom[2697] = 'b001101010;assign rom[2698] = 'b001011000;assign rom[2699] = 'b101001000;assign rom[2700] = 'b000101011;assign rom[2701] = 'b110000010;assign rom[2702] = 'b111000000;assign rom[2703] = 'b101001100;assign rom[2704] = 'b001001010;assign rom[2705] = 'b111111000;assign rom[2706] = 'b111101000;assign rom[2707] = 'b101001111;assign rom[2708] = 'b000111010;assign rom[2709] = 'b101110110;assign rom[2710] = 'b101100010;assign rom[2711] = 'b101001100;assign rom[2712] = 'b001001010;assign rom[2713] = 'b111011010;assign rom[2714] = 'b111011010;assign rom[2715] = 'b111011010;assign rom[2716] = 'b111011010;assign rom[2717] = 'b111011000;assign rom[2718] = 'b111011000;assign rom[2719] = 'b111011000;assign rom[2720] = 'b111011000;assign rom[2721] = 'b101111000;assign rom[2722] = 'b000110011;assign rom[2723] = 'b110000010;assign rom[2724] = 'b001101010;assign rom[2725] = 'b001011000;assign rom[2726] = 'b101001000;assign rom[2727] = 'b000101011;assign rom[2728] = 'b110000010;assign rom[2729] = 'b111000000;assign rom[2730] = 'b101001100;assign rom[2731] = 'b001001010;assign rom[2732] = 'b111111000;assign rom[2733] = 'b111101000;assign rom[2734] = 'b101001111;assign rom[2735] = 'b000111010;assign rom[2736] = 'b101110110;assign rom[2737] = 'b101100010;assign rom[2738] = 'b101001100;assign rom[2739] = 'b001001010;assign rom[2740] = 'b111011010;assign rom[2741] = 'b111011010;assign rom[2742] = 'b111011010;assign rom[2743] = 'b111011010;assign rom[2744] = 'b111011000;assign rom[2745] = 'b111011000;assign rom[2746] = 'b111011000;assign rom[2747] = 'b111011000;assign rom[2748] = 'b101111000;assign rom[2749] = 'b000110011;assign rom[2750] = 'b110000010;assign rom[2751] = 'b001101010;assign rom[2752] = 'b001011000;assign rom[2753] = 'b101001000;assign rom[2754] = 'b000101011;assign rom[2755] = 'b110000010;assign rom[2756] = 'b111000000;assign rom[2757] = 'b101001100;assign rom[2758] = 'b001001010;assign rom[2759] = 'b111111000;assign rom[2760] = 'b111101000;assign rom[2761] = 'b101001111;assign rom[2762] = 'b000111010;assign rom[2763] = 'b101110110;assign rom[2764] = 'b101100010;assign rom[2765] = 'b101001100;assign rom[2766] = 'b001001010;assign rom[2767] = 'b111011010;assign rom[2768] = 'b111011010;assign rom[2769] = 'b111011010;assign rom[2770] = 'b111011010;assign rom[2771] = 'b111011000;assign rom[2772] = 'b111011000;assign rom[2773] = 'b111011000;assign rom[2774] = 'b111011000;assign rom[2775] = 'b101111000;assign rom[2776] = 'b000110011;assign rom[2777] = 'b110000010;assign rom[2778] = 'b001101010;assign rom[2779] = 'b001011000;assign rom[2780] = 'b101001000;assign rom[2781] = 'b000101011;assign rom[2782] = 'b110000010;assign rom[2783] = 'b111000000;assign rom[2784] = 'b101001100;assign rom[2785] = 'b001001010;assign rom[2786] = 'b111111000;assign rom[2787] = 'b111101000;assign rom[2788] = 'b101001111;assign rom[2789] = 'b000111010;assign rom[2790] = 'b101110110;assign rom[2791] = 'b101100010;assign rom[2792] = 'b101001100;assign rom[2793] = 'b001001010;assign rom[2794] = 'b111011010;assign rom[2795] = 'b111011010;assign rom[2796] = 'b111011010;assign rom[2797] = 'b111011010;assign rom[2798] = 'b111011000;assign rom[2799] = 'b111011000;assign rom[2800] = 'b111011000;assign rom[2801] = 'b111011000;assign rom[2802] = 'b101111000;assign rom[2803] = 'b000110011;assign rom[2804] = 'b110000010;assign rom[2805] = 'b001101010;assign rom[2806] = 'b001011000;assign rom[2807] = 'b101001000;assign rom[2808] = 'b000101011;assign rom[2809] = 'b110000010;assign rom[2810] = 'b111000000;assign rom[2811] = 'b101001100;assign rom[2812] = 'b001001010;assign rom[2813] = 'b111111000;assign rom[2814] = 'b111101000;assign rom[2815] = 'b101001111;assign rom[2816] = 'b000111010;assign rom[2817] = 'b101110110;assign rom[2818] = 'b101100010;assign rom[2819] = 'b101001100;assign rom[2820] = 'b001001010;assign rom[2821] = 'b111011010;assign rom[2822] = 'b111011010;assign rom[2823] = 'b111011010;assign rom[2824] = 'b111011010;assign rom[2825] = 'b111011000;assign rom[2826] = 'b111011000;assign rom[2827] = 'b111011000;assign rom[2828] = 'b111011000;assign rom[2829] = 'b101111000;assign rom[2830] = 'b000110011;assign rom[2831] = 'b110000010;assign rom[2832] = 'b001101010;assign rom[2833] = 'b001011000;assign rom[2834] = 'b101001000;assign rom[2835] = 'b000101011;assign rom[2836] = 'b110000010;assign rom[2837] = 'b111000000;assign rom[2838] = 'b101001100;assign rom[2839] = 'b001001010;assign rom[2840] = 'b111111000;assign rom[2841] = 'b111101000;assign rom[2842] = 'b101001111;assign rom[2843] = 'b000111010;assign rom[2844] = 'b101110110;assign rom[2845] = 'b101100010;assign rom[2846] = 'b101001100;assign rom[2847] = 'b001001010;assign rom[2848] = 'b111011010;assign rom[2849] = 'b111011010;assign rom[2850] = 'b111011010;assign rom[2851] = 'b111011010;assign rom[2852] = 'b111011000;assign rom[2853] = 'b111011000;assign rom[2854] = 'b111011000;assign rom[2855] = 'b111011000;assign rom[2856] = 'b101111000;assign rom[2857] = 'b000110011;assign rom[2858] = 'b110000010;assign rom[2859] = 'b001101010;assign rom[2860] = 'b001011000;assign rom[2861] = 'b101001000;assign rom[2862] = 'b000101011;assign rom[2863] = 'b110000010;assign rom[2864] = 'b111000000;assign rom[2865] = 'b101001100;assign rom[2866] = 'b001001010;assign rom[2867] = 'b111111000;assign rom[2868] = 'b111101000;assign rom[2869] = 'b101001111;assign rom[2870] = 'b000111010;assign rom[2871] = 'b101110110;assign rom[2872] = 'b101100010;assign rom[2873] = 'b101001100;assign rom[2874] = 'b001001010;assign rom[2875] = 'b111011010;assign rom[2876] = 'b111011010;assign rom[2877] = 'b111011010;assign rom[2878] = 'b111011010;assign rom[2879] = 'b111011000;assign rom[2880] = 'b111011000;assign rom[2881] = 'b111011000;assign rom[2882] = 'b111011000;assign rom[2883] = 'b101111000;assign rom[2884] = 'b000110011;assign rom[2885] = 'b110000010;assign rom[2886] = 'b001101010;assign rom[2887] = 'b001011000;assign rom[2888] = 'b101001000;assign rom[2889] = 'b000101011;assign rom[2890] = 'b110000010;assign rom[2891] = 'b111000000;assign rom[2892] = 'b101001100;assign rom[2893] = 'b001001010;assign rom[2894] = 'b111111000;assign rom[2895] = 'b111101000;assign rom[2896] = 'b101001111;assign rom[2897] = 'b000111010;assign rom[2898] = 'b101110110;assign rom[2899] = 'b101100010;assign rom[2900] = 'b101001100;assign rom[2901] = 'b001001010;assign rom[2902] = 'b111011010;assign rom[2903] = 'b111011010;assign rom[2904] = 'b111011010;assign rom[2905] = 'b111011010;assign rom[2906] = 'b111011000;assign rom[2907] = 'b111011000;assign rom[2908] = 'b111011000;assign rom[2909] = 'b111011000;assign rom[2910] = 'b101111000;assign rom[2911] = 'b000110011;assign rom[2912] = 'b110000010;assign rom[2913] = 'b001101010;assign rom[2914] = 'b001011000;assign rom[2915] = 'b101001000;assign rom[2916] = 'b000101011;assign rom[2917] = 'b110000010;assign rom[2918] = 'b111000000;assign rom[2919] = 'b101001100;assign rom[2920] = 'b001001010;assign rom[2921] = 'b001000110;assign rom[2922] = 'b001100100;assign rom[2923] = 'b101100010;assign rom[2924] = 'b101001100;assign rom[2925] = 'b001001010;assign rom[2926] = 'b111011010;assign rom[2927] = 'b111011010;assign rom[2928] = 'b111011010;assign rom[2929] = 'b111011010;assign rom[2930] = 'b111011000;assign rom[2931] = 'b111011000;assign rom[2932] = 'b111011000;assign rom[2933] = 'b111011000;assign rom[2934] = 'b101111000;assign rom[2935] = 'b000110011;assign rom[2936] = 'b110000010;assign rom[2937] = 'b001101010;assign rom[2938] = 'b001011000;assign rom[2939] = 'b101001000;assign rom[2940] = 'b000101011;assign rom[2941] = 'b110000010;assign rom[2942] = 'b111000000;assign rom[2943] = 'b101001100;assign rom[2944] = 'b001001010;assign rom[2945] = 'b111111000;assign rom[2946] = 'b111101000;assign rom[2947] = 'b101001111;assign rom[2948] = 'b000111010;assign rom[2949] = 'b101110110;assign rom[2950] = 'b101100010;assign rom[2951] = 'b101001100;assign rom[2952] = 'b001001010;assign rom[2953] = 'b111011010;assign rom[2954] = 'b111011010;assign rom[2955] = 'b111011010;assign rom[2956] = 'b111011010;assign rom[2957] = 'b111011000;assign rom[2958] = 'b111011000;assign rom[2959] = 'b111011000;assign rom[2960] = 'b111011000;assign rom[2961] = 'b101111000;assign rom[2962] = 'b000110011;assign rom[2963] = 'b110000010;assign rom[2964] = 'b001101010;assign rom[2965] = 'b001011000;assign rom[2966] = 'b101001000;assign rom[2967] = 'b000101011;assign rom[2968] = 'b110000010;assign rom[2969] = 'b111000000;assign rom[2970] = 'b101001100;assign rom[2971] = 'b001001010;assign rom[2972] = 'b111111000;assign rom[2973] = 'b111101000;assign rom[2974] = 'b101001111;assign rom[2975] = 'b000111010;assign rom[2976] = 'b101110110;assign rom[2977] = 'b101100010;assign rom[2978] = 'b101001100;assign rom[2979] = 'b001001010;assign rom[2980] = 'b111011010;assign rom[2981] = 'b111011010;assign rom[2982] = 'b111011010;assign rom[2983] = 'b111011010;assign rom[2984] = 'b111011000;assign rom[2985] = 'b111011000;assign rom[2986] = 'b111011000;assign rom[2987] = 'b111011000;assign rom[2988] = 'b101111000;assign rom[2989] = 'b000110011;assign rom[2990] = 'b110000010;assign rom[2991] = 'b001101010;assign rom[2992] = 'b001011000;assign rom[2993] = 'b101001000;assign rom[2994] = 'b000101011;assign rom[2995] = 'b110000010;assign rom[2996] = 'b111000000;assign rom[2997] = 'b101001100;assign rom[2998] = 'b001001010;assign rom[2999] = 'b111111000;assign rom[3000] = 'b111101000;assign rom[3001] = 'b101001111;assign rom[3002] = 'b000111010;assign rom[3003] = 'b101110110;assign rom[3004] = 'b101100010;assign rom[3005] = 'b101001100;assign rom[3006] = 'b001001010;assign rom[3007] = 'b111011010;assign rom[3008] = 'b111011010;assign rom[3009] = 'b111011010;assign rom[3010] = 'b111011010;assign rom[3011] = 'b111011000;assign rom[3012] = 'b111011000;assign rom[3013] = 'b111011000;assign rom[3014] = 'b111011000;assign rom[3015] = 'b101111000;assign rom[3016] = 'b000110011;assign rom[3017] = 'b110000010;assign rom[3018] = 'b001101010;assign rom[3019] = 'b001011000;assign rom[3020] = 'b101001000;assign rom[3021] = 'b000101011;assign rom[3022] = 'b110000010;assign rom[3023] = 'b111000000;assign rom[3024] = 'b101001100;assign rom[3025] = 'b001001010;assign rom[3026] = 'b111111000;assign rom[3027] = 'b111101000;assign rom[3028] = 'b101001111;assign rom[3029] = 'b000111010;assign rom[3030] = 'b101110110;assign rom[3031] = 'b101100010;assign rom[3032] = 'b101001100;assign rom[3033] = 'b001001010;assign rom[3034] = 'b111011010;assign rom[3035] = 'b111011010;assign rom[3036] = 'b111011010;assign rom[3037] = 'b111011010;assign rom[3038] = 'b111011000;assign rom[3039] = 'b111011000;assign rom[3040] = 'b111011000;assign rom[3041] = 'b111011000;assign rom[3042] = 'b101111000;assign rom[3043] = 'b000110011;assign rom[3044] = 'b110000010;assign rom[3045] = 'b001101010;assign rom[3046] = 'b001011000;assign rom[3047] = 'b101001000;assign rom[3048] = 'b000101011;assign rom[3049] = 'b110000010;assign rom[3050] = 'b111000000;assign rom[3051] = 'b101001100;assign rom[3052] = 'b001001010;assign rom[3053] = 'b111111000;assign rom[3054] = 'b111101000;assign rom[3055] = 'b101001111;assign rom[3056] = 'b000111010;assign rom[3057] = 'b101110110;assign rom[3058] = 'b101100010;assign rom[3059] = 'b101001100;assign rom[3060] = 'b001001010;assign rom[3061] = 'b111011010;assign rom[3062] = 'b111011010;assign rom[3063] = 'b111011010;assign rom[3064] = 'b111011010;assign rom[3065] = 'b111011000;assign rom[3066] = 'b111011000;assign rom[3067] = 'b111011000;assign rom[3068] = 'b111011000;assign rom[3069] = 'b101111000;assign rom[3070] = 'b000110011;assign rom[3071] = 'b110000010;assign rom[3072] = 'b001101010;assign rom[3073] = 'b001011000;assign rom[3074] = 'b101001000;assign rom[3075] = 'b000101011;assign rom[3076] = 'b110000010;assign rom[3077] = 'b111000000;assign rom[3078] = 'b101001100;assign rom[3079] = 'b001001010;assign rom[3080] = 'b111111000;assign rom[3081] = 'b111101000;assign rom[3082] = 'b101001111;assign rom[3083] = 'b000111010;assign rom[3084] = 'b101110110;assign rom[3085] = 'b101100010;assign rom[3086] = 'b101001100;assign rom[3087] = 'b001001010;assign rom[3088] = 'b111011010;assign rom[3089] = 'b111011010;assign rom[3090] = 'b111011010;assign rom[3091] = 'b111011010;assign rom[3092] = 'b111011000;assign rom[3093] = 'b111011000;assign rom[3094] = 'b111011000;assign rom[3095] = 'b111011000;assign rom[3096] = 'b101111000;assign rom[3097] = 'b000110011;assign rom[3098] = 'b110000010;assign rom[3099] = 'b001101010;assign rom[3100] = 'b001011000;assign rom[3101] = 'b101001000;assign rom[3102] = 'b000101011;assign rom[3103] = 'b110000010;assign rom[3104] = 'b111000000;assign rom[3105] = 'b101001100;assign rom[3106] = 'b001001010;assign rom[3107] = 'b111111000;assign rom[3108] = 'b111101000;assign rom[3109] = 'b101001111;assign rom[3110] = 'b000111010;assign rom[3111] = 'b101110110;assign rom[3112] = 'b101100010;assign rom[3113] = 'b101001100;assign rom[3114] = 'b001001010;assign rom[3115] = 'b111011010;assign rom[3116] = 'b111011010;assign rom[3117] = 'b111011010;assign rom[3118] = 'b111011010;assign rom[3119] = 'b111011000;assign rom[3120] = 'b111011000;assign rom[3121] = 'b111011000;assign rom[3122] = 'b111011000;assign rom[3123] = 'b101111000;assign rom[3124] = 'b000110011;assign rom[3125] = 'b110000010;assign rom[3126] = 'b001101010;assign rom[3127] = 'b001011000;assign rom[3128] = 'b101001000;assign rom[3129] = 'b000101011;assign rom[3130] = 'b110000010;assign rom[3131] = 'b111000000;assign rom[3132] = 'b101001100;assign rom[3133] = 'b001001010;assign rom[3134] = 'b111111000;assign rom[3135] = 'b111101000;assign rom[3136] = 'b101001111;assign rom[3137] = 'b000111010;assign rom[3138] = 'b101110110;assign rom[3139] = 'b101100010;assign rom[3140] = 'b101001100;assign rom[3141] = 'b001001010;assign rom[3142] = 'b111011010;assign rom[3143] = 'b111011010;assign rom[3144] = 'b111011010;assign rom[3145] = 'b111011010;assign rom[3146] = 'b111011000;assign rom[3147] = 'b111011000;assign rom[3148] = 'b111011000;assign rom[3149] = 'b111011000;assign rom[3150] = 'b101111000;assign rom[3151] = 'b000110011;assign rom[3152] = 'b110000010;assign rom[3153] = 'b001101010;assign rom[3154] = 'b001011000;assign rom[3155] = 'b101001000;assign rom[3156] = 'b000101011;assign rom[3157] = 'b110000010;assign rom[3158] = 'b111000000;assign rom[3159] = 'b101001100;assign rom[3160] = 'b001001010;assign rom[3161] = 'b001000110;assign rom[3162] = 'b001100100;assign rom[3163] = 'b101100010;assign rom[3164] = 'b101001100;assign rom[3165] = 'b001001010;assign rom[3166] = 'b111011010;assign rom[3167] = 'b111011010;assign rom[3168] = 'b111011010;assign rom[3169] = 'b111011010;assign rom[3170] = 'b111011000;assign rom[3171] = 'b111011000;assign rom[3172] = 'b111011000;assign rom[3173] = 'b111011000;assign rom[3174] = 'b101111000;assign rom[3175] = 'b000110011;assign rom[3176] = 'b110000010;assign rom[3177] = 'b001101010;assign rom[3178] = 'b001011000;assign rom[3179] = 'b101001000;assign rom[3180] = 'b000101011;assign rom[3181] = 'b110000010;assign rom[3182] = 'b111000000;assign rom[3183] = 'b101001100;assign rom[3184] = 'b001001010;assign rom[3185] = 'b111111000;assign rom[3186] = 'b111101000;assign rom[3187] = 'b101001111;assign rom[3188] = 'b000111010;assign rom[3189] = 'b101110110;assign rom[3190] = 'b101100010;assign rom[3191] = 'b101001100;assign rom[3192] = 'b001001010;assign rom[3193] = 'b111011010;assign rom[3194] = 'b111011010;assign rom[3195] = 'b111011010;assign rom[3196] = 'b111011010;assign rom[3197] = 'b111011000;assign rom[3198] = 'b111011000;assign rom[3199] = 'b111011000;assign rom[3200] = 'b111011000;assign rom[3201] = 'b101111000;assign rom[3202] = 'b000110011;assign rom[3203] = 'b110000010;assign rom[3204] = 'b001101010;assign rom[3205] = 'b001011000;assign rom[3206] = 'b101001000;assign rom[3207] = 'b000101011;assign rom[3208] = 'b110000010;assign rom[3209] = 'b111000000;assign rom[3210] = 'b101001100;assign rom[3211] = 'b001001010;assign rom[3212] = 'b111111000;assign rom[3213] = 'b111101000;assign rom[3214] = 'b101001111;assign rom[3215] = 'b000111010;assign rom[3216] = 'b101110110;assign rom[3217] = 'b101100010;assign rom[3218] = 'b101001100;assign rom[3219] = 'b001001010;assign rom[3220] = 'b111011010;assign rom[3221] = 'b111011010;assign rom[3222] = 'b111011010;assign rom[3223] = 'b111011010;assign rom[3224] = 'b111011000;assign rom[3225] = 'b111011000;assign rom[3226] = 'b111011000;assign rom[3227] = 'b111011000;assign rom[3228] = 'b101111000;assign rom[3229] = 'b000110011;assign rom[3230] = 'b110000010;assign rom[3231] = 'b001101010;assign rom[3232] = 'b001011000;assign rom[3233] = 'b101001000;assign rom[3234] = 'b000101011;assign rom[3235] = 'b110000010;assign rom[3236] = 'b111000000;assign rom[3237] = 'b101001100;assign rom[3238] = 'b001001010;assign rom[3239] = 'b111111000;assign rom[3240] = 'b111101000;assign rom[3241] = 'b101001111;assign rom[3242] = 'b000111010;assign rom[3243] = 'b101110110;assign rom[3244] = 'b101100010;assign rom[3245] = 'b101001100;assign rom[3246] = 'b001001010;assign rom[3247] = 'b111011010;assign rom[3248] = 'b111011010;assign rom[3249] = 'b111011010;assign rom[3250] = 'b111011010;assign rom[3251] = 'b111011000;assign rom[3252] = 'b111011000;assign rom[3253] = 'b111011000;assign rom[3254] = 'b111011000;assign rom[3255] = 'b101111000;assign rom[3256] = 'b000110011;assign rom[3257] = 'b110000010;assign rom[3258] = 'b001101010;assign rom[3259] = 'b001011000;assign rom[3260] = 'b101001000;assign rom[3261] = 'b000101011;assign rom[3262] = 'b110000010;assign rom[3263] = 'b111000000;assign rom[3264] = 'b101001100;assign rom[3265] = 'b001001010;assign rom[3266] = 'b111111000;assign rom[3267] = 'b111101000;assign rom[3268] = 'b101001111;assign rom[3269] = 'b000111010;assign rom[3270] = 'b101110110;assign rom[3271] = 'b101100010;assign rom[3272] = 'b101001100;assign rom[3273] = 'b001001010;assign rom[3274] = 'b111011010;assign rom[3275] = 'b111011010;assign rom[3276] = 'b111011010;assign rom[3277] = 'b111011010;assign rom[3278] = 'b111011000;assign rom[3279] = 'b111011000;assign rom[3280] = 'b111011000;assign rom[3281] = 'b111011000;assign rom[3282] = 'b101111000;assign rom[3283] = 'b000110011;assign rom[3284] = 'b110000010;assign rom[3285] = 'b001101010;assign rom[3286] = 'b001011000;assign rom[3287] = 'b101001000;assign rom[3288] = 'b000101011;assign rom[3289] = 'b110000010;assign rom[3290] = 'b111000000;assign rom[3291] = 'b101001100;assign rom[3292] = 'b001001010;assign rom[3293] = 'b111111000;assign rom[3294] = 'b111101000;assign rom[3295] = 'b101001111;assign rom[3296] = 'b000111010;assign rom[3297] = 'b101110110;assign rom[3298] = 'b101100010;assign rom[3299] = 'b101001100;assign rom[3300] = 'b001001010;assign rom[3301] = 'b111011010;assign rom[3302] = 'b111011010;assign rom[3303] = 'b111011010;assign rom[3304] = 'b111011010;assign rom[3305] = 'b111011000;assign rom[3306] = 'b111011000;assign rom[3307] = 'b111011000;assign rom[3308] = 'b111011000;assign rom[3309] = 'b101111000;assign rom[3310] = 'b000110011;assign rom[3311] = 'b110000010;assign rom[3312] = 'b001101010;assign rom[3313] = 'b001011000;assign rom[3314] = 'b101001000;assign rom[3315] = 'b000101011;assign rom[3316] = 'b110000010;assign rom[3317] = 'b111000000;assign rom[3318] = 'b101001100;assign rom[3319] = 'b001001010;assign rom[3320] = 'b111111000;assign rom[3321] = 'b111101000;assign rom[3322] = 'b101001111;assign rom[3323] = 'b000111010;assign rom[3324] = 'b101110110;assign rom[3325] = 'b101100010;assign rom[3326] = 'b101001100;assign rom[3327] = 'b001001010;assign rom[3328] = 'b111011010;assign rom[3329] = 'b111011010;assign rom[3330] = 'b111011010;assign rom[3331] = 'b111011010;assign rom[3332] = 'b111011000;assign rom[3333] = 'b111011000;assign rom[3334] = 'b111011000;assign rom[3335] = 'b111011000;assign rom[3336] = 'b101111000;assign rom[3337] = 'b000110011;assign rom[3338] = 'b110000010;assign rom[3339] = 'b001101010;assign rom[3340] = 'b001011000;assign rom[3341] = 'b101001000;assign rom[3342] = 'b000101011;assign rom[3343] = 'b110000010;assign rom[3344] = 'b111000000;assign rom[3345] = 'b101001100;assign rom[3346] = 'b001001010;assign rom[3347] = 'b111111000;assign rom[3348] = 'b111101000;assign rom[3349] = 'b101001111;assign rom[3350] = 'b000111010;assign rom[3351] = 'b101110110;assign rom[3352] = 'b101100010;assign rom[3353] = 'b101001100;assign rom[3354] = 'b001001010;assign rom[3355] = 'b111011010;assign rom[3356] = 'b111011010;assign rom[3357] = 'b111011010;assign rom[3358] = 'b111011010;assign rom[3359] = 'b111011000;assign rom[3360] = 'b111011000;assign rom[3361] = 'b111011000;assign rom[3362] = 'b111011000;assign rom[3363] = 'b101111000;assign rom[3364] = 'b000110011;assign rom[3365] = 'b110000010;assign rom[3366] = 'b001101010;assign rom[3367] = 'b001011000;assign rom[3368] = 'b101001000;assign rom[3369] = 'b000101011;assign rom[3370] = 'b110000010;assign rom[3371] = 'b111000000;assign rom[3372] = 'b101001100;assign rom[3373] = 'b001001010;assign rom[3374] = 'b111111000;assign rom[3375] = 'b111101000;assign rom[3376] = 'b101001111;assign rom[3377] = 'b000111010;assign rom[3378] = 'b101110110;assign rom[3379] = 'b101100010;assign rom[3380] = 'b101001100;assign rom[3381] = 'b001001010;assign rom[3382] = 'b111011010;assign rom[3383] = 'b111011010;assign rom[3384] = 'b111011010;assign rom[3385] = 'b111011010;assign rom[3386] = 'b111011000;assign rom[3387] = 'b111011000;assign rom[3388] = 'b111011000;assign rom[3389] = 'b111011000;assign rom[3390] = 'b101111000;assign rom[3391] = 'b000110011;assign rom[3392] = 'b110000010;assign rom[3393] = 'b001101010;assign rom[3394] = 'b001011000;assign rom[3395] = 'b101001000;assign rom[3396] = 'b000101011;assign rom[3397] = 'b110000010;assign rom[3398] = 'b111000000;assign rom[3399] = 'b101001100;assign rom[3400] = 'b001001010;assign rom[3401] = 'b001000110;assign rom[3402] = 'b001100100;assign rom[3403] = 'b101100010;assign rom[3404] = 'b101001100;assign rom[3405] = 'b001001010;assign rom[3406] = 'b111011010;assign rom[3407] = 'b111011010;assign rom[3408] = 'b111011010;assign rom[3409] = 'b111011010;assign rom[3410] = 'b111011000;assign rom[3411] = 'b111011000;assign rom[3412] = 'b111011000;assign rom[3413] = 'b111011000;assign rom[3414] = 'b101111000;assign rom[3415] = 'b000110011;assign rom[3416] = 'b110000010;assign rom[3417] = 'b001101010;assign rom[3418] = 'b001011000;assign rom[3419] = 'b101001000;assign rom[3420] = 'b000101011;assign rom[3421] = 'b110000010;assign rom[3422] = 'b111000000;assign rom[3423] = 'b101001100;assign rom[3424] = 'b001001010;assign rom[3425] = 'b111111000;assign rom[3426] = 'b111101000;assign rom[3427] = 'b101001111;assign rom[3428] = 'b000111010;assign rom[3429] = 'b101110110;assign rom[3430] = 'b101100010;assign rom[3431] = 'b101001100;assign rom[3432] = 'b001001010;assign rom[3433] = 'b111011010;assign rom[3434] = 'b111011010;assign rom[3435] = 'b111011010;assign rom[3436] = 'b111011010;assign rom[3437] = 'b111011000;assign rom[3438] = 'b111011000;assign rom[3439] = 'b111011000;assign rom[3440] = 'b111011000;assign rom[3441] = 'b101111000;assign rom[3442] = 'b000110011;assign rom[3443] = 'b110000010;assign rom[3444] = 'b001101010;assign rom[3445] = 'b001011000;assign rom[3446] = 'b101001000;assign rom[3447] = 'b000101011;assign rom[3448] = 'b110000010;assign rom[3449] = 'b111000000;assign rom[3450] = 'b101001100;assign rom[3451] = 'b001001010;assign rom[3452] = 'b111111000;assign rom[3453] = 'b111101000;assign rom[3454] = 'b101001111;assign rom[3455] = 'b000111010;assign rom[3456] = 'b101110110;assign rom[3457] = 'b101100010;assign rom[3458] = 'b101001100;assign rom[3459] = 'b001001010;assign rom[3460] = 'b111011010;assign rom[3461] = 'b111011010;assign rom[3462] = 'b111011010;assign rom[3463] = 'b111011010;assign rom[3464] = 'b111011000;assign rom[3465] = 'b111011000;assign rom[3466] = 'b111011000;assign rom[3467] = 'b111011000;assign rom[3468] = 'b101111000;assign rom[3469] = 'b000110011;assign rom[3470] = 'b110000010;assign rom[3471] = 'b001101010;assign rom[3472] = 'b001011000;assign rom[3473] = 'b101001000;assign rom[3474] = 'b000101011;assign rom[3475] = 'b110000010;assign rom[3476] = 'b111000000;assign rom[3477] = 'b101001100;assign rom[3478] = 'b001001010;assign rom[3479] = 'b111111000;assign rom[3480] = 'b111101000;assign rom[3481] = 'b101001111;assign rom[3482] = 'b000111010;assign rom[3483] = 'b101110110;assign rom[3484] = 'b101100010;assign rom[3485] = 'b101001100;assign rom[3486] = 'b001001010;assign rom[3487] = 'b111011010;assign rom[3488] = 'b111011010;assign rom[3489] = 'b111011010;assign rom[3490] = 'b111011010;assign rom[3491] = 'b111011000;assign rom[3492] = 'b111011000;assign rom[3493] = 'b111011000;assign rom[3494] = 'b111011000;assign rom[3495] = 'b101111000;assign rom[3496] = 'b000110011;assign rom[3497] = 'b110000010;assign rom[3498] = 'b001101010;assign rom[3499] = 'b001011000;assign rom[3500] = 'b101001000;assign rom[3501] = 'b000101011;assign rom[3502] = 'b110000010;assign rom[3503] = 'b111000000;assign rom[3504] = 'b101001100;assign rom[3505] = 'b001001010;assign rom[3506] = 'b111111000;assign rom[3507] = 'b111101000;assign rom[3508] = 'b101001111;assign rom[3509] = 'b000111010;assign rom[3510] = 'b101110110;assign rom[3511] = 'b101100010;assign rom[3512] = 'b101001100;assign rom[3513] = 'b001001010;assign rom[3514] = 'b111011010;assign rom[3515] = 'b111011010;assign rom[3516] = 'b111011010;assign rom[3517] = 'b111011010;assign rom[3518] = 'b111011000;assign rom[3519] = 'b111011000;assign rom[3520] = 'b111011000;assign rom[3521] = 'b111011000;assign rom[3522] = 'b101111000;assign rom[3523] = 'b000110011;assign rom[3524] = 'b110000010;assign rom[3525] = 'b001101010;assign rom[3526] = 'b001011000;assign rom[3527] = 'b101001000;assign rom[3528] = 'b000101011;assign rom[3529] = 'b110000010;assign rom[3530] = 'b111000000;assign rom[3531] = 'b101001100;assign rom[3532] = 'b001001010;assign rom[3533] = 'b111111000;assign rom[3534] = 'b111101000;assign rom[3535] = 'b101001111;assign rom[3536] = 'b000111010;assign rom[3537] = 'b101110110;assign rom[3538] = 'b101100010;assign rom[3539] = 'b101001100;assign rom[3540] = 'b001001010;assign rom[3541] = 'b111011010;assign rom[3542] = 'b111011010;assign rom[3543] = 'b111011010;assign rom[3544] = 'b111011010;assign rom[3545] = 'b111011000;assign rom[3546] = 'b111011000;assign rom[3547] = 'b111011000;assign rom[3548] = 'b111011000;assign rom[3549] = 'b101111000;assign rom[3550] = 'b000110011;assign rom[3551] = 'b110000010;assign rom[3552] = 'b001101010;assign rom[3553] = 'b001011000;assign rom[3554] = 'b101001000;assign rom[3555] = 'b000101011;assign rom[3556] = 'b110000010;assign rom[3557] = 'b111000000;assign rom[3558] = 'b101001100;assign rom[3559] = 'b001001010;assign rom[3560] = 'b111111000;assign rom[3561] = 'b111101000;assign rom[3562] = 'b101001111;assign rom[3563] = 'b000111010;assign rom[3564] = 'b101110110;assign rom[3565] = 'b101100010;assign rom[3566] = 'b101001100;assign rom[3567] = 'b001001010;assign rom[3568] = 'b111011010;assign rom[3569] = 'b111011010;assign rom[3570] = 'b111011010;assign rom[3571] = 'b111011010;assign rom[3572] = 'b111011000;assign rom[3573] = 'b111011000;assign rom[3574] = 'b111011000;assign rom[3575] = 'b111011000;assign rom[3576] = 'b101111000;assign rom[3577] = 'b000110011;assign rom[3578] = 'b110000010;assign rom[3579] = 'b001101010;assign rom[3580] = 'b001011000;assign rom[3581] = 'b101001000;assign rom[3582] = 'b000101011;assign rom[3583] = 'b110000010;assign rom[3584] = 'b111000000;assign rom[3585] = 'b101001100;assign rom[3586] = 'b001001010;assign rom[3587] = 'b111111000;assign rom[3588] = 'b111101000;assign rom[3589] = 'b101001111;assign rom[3590] = 'b000111010;assign rom[3591] = 'b101110110;assign rom[3592] = 'b101100010;assign rom[3593] = 'b101001100;assign rom[3594] = 'b001001010;assign rom[3595] = 'b111011010;assign rom[3596] = 'b111011010;assign rom[3597] = 'b111011010;assign rom[3598] = 'b111011010;assign rom[3599] = 'b111011000;assign rom[3600] = 'b111011000;assign rom[3601] = 'b111011000;assign rom[3602] = 'b111011000;assign rom[3603] = 'b101111000;assign rom[3604] = 'b000110011;assign rom[3605] = 'b110000010;assign rom[3606] = 'b001101010;assign rom[3607] = 'b001011000;assign rom[3608] = 'b101001000;assign rom[3609] = 'b000101011;assign rom[3610] = 'b110000010;assign rom[3611] = 'b111000000;assign rom[3612] = 'b101001100;assign rom[3613] = 'b001001010;assign rom[3614] = 'b111111000;assign rom[3615] = 'b111101000;assign rom[3616] = 'b101001111;assign rom[3617] = 'b000111010;assign rom[3618] = 'b101110110;assign rom[3619] = 'b101100010;assign rom[3620] = 'b101001100;assign rom[3621] = 'b001001010;assign rom[3622] = 'b111011010;assign rom[3623] = 'b111011010;assign rom[3624] = 'b111011010;assign rom[3625] = 'b111011010;assign rom[3626] = 'b111011000;assign rom[3627] = 'b111011000;assign rom[3628] = 'b111011000;assign rom[3629] = 'b111011000;assign rom[3630] = 'b101111000;assign rom[3631] = 'b000110011;assign rom[3632] = 'b110000010;assign rom[3633] = 'b001101010;assign rom[3634] = 'b001011000;assign rom[3635] = 'b101001000;assign rom[3636] = 'b000101011;assign rom[3637] = 'b110000010;assign rom[3638] = 'b111000000;assign rom[3639] = 'b101001100;assign rom[3640] = 'b001001010;assign rom[3641] = 'b001000110;assign rom[3642] = 'b001100100;assign rom[3643] = 'b101100010;assign rom[3644] = 'b101001100;assign rom[3645] = 'b001001010;assign rom[3646] = 'b111011010;assign rom[3647] = 'b111011010;assign rom[3648] = 'b111011010;assign rom[3649] = 'b111011010;assign rom[3650] = 'b111011000;assign rom[3651] = 'b111011000;assign rom[3652] = 'b111011000;assign rom[3653] = 'b111011000;assign rom[3654] = 'b101111000;assign rom[3655] = 'b000110011;assign rom[3656] = 'b110000010;assign rom[3657] = 'b001101010;assign rom[3658] = 'b001011000;assign rom[3659] = 'b101001000;assign rom[3660] = 'b000101011;assign rom[3661] = 'b110000010;assign rom[3662] = 'b111000000;assign rom[3663] = 'b101001100;assign rom[3664] = 'b001001010;assign rom[3665] = 'b111111000;assign rom[3666] = 'b111101000;assign rom[3667] = 'b101001111;assign rom[3668] = 'b000111010;assign rom[3669] = 'b101110110;assign rom[3670] = 'b101100010;assign rom[3671] = 'b101001100;assign rom[3672] = 'b001001010;assign rom[3673] = 'b111011010;assign rom[3674] = 'b111011010;assign rom[3675] = 'b111011010;assign rom[3676] = 'b111011010;assign rom[3677] = 'b111011000;assign rom[3678] = 'b111011000;assign rom[3679] = 'b111011000;assign rom[3680] = 'b111011000;assign rom[3681] = 'b101111000;assign rom[3682] = 'b000110011;assign rom[3683] = 'b110000010;assign rom[3684] = 'b001101010;assign rom[3685] = 'b001011000;assign rom[3686] = 'b101001000;assign rom[3687] = 'b000101011;assign rom[3688] = 'b110000010;assign rom[3689] = 'b111000000;assign rom[3690] = 'b101001100;assign rom[3691] = 'b001001010;assign rom[3692] = 'b111111000;assign rom[3693] = 'b111101000;assign rom[3694] = 'b101001111;assign rom[3695] = 'b000111010;assign rom[3696] = 'b101110110;assign rom[3697] = 'b101100010;assign rom[3698] = 'b101001100;assign rom[3699] = 'b001001010;assign rom[3700] = 'b111011010;assign rom[3701] = 'b111011010;assign rom[3702] = 'b111011010;assign rom[3703] = 'b111011010;assign rom[3704] = 'b111011000;assign rom[3705] = 'b111011000;assign rom[3706] = 'b111011000;assign rom[3707] = 'b111011000;assign rom[3708] = 'b101111000;assign rom[3709] = 'b000110011;assign rom[3710] = 'b110000010;assign rom[3711] = 'b001101010;assign rom[3712] = 'b001011000;assign rom[3713] = 'b101001000;assign rom[3714] = 'b000101011;assign rom[3715] = 'b110000010;assign rom[3716] = 'b111000000;assign rom[3717] = 'b101001100;assign rom[3718] = 'b001001010;assign rom[3719] = 'b111111000;assign rom[3720] = 'b111101000;assign rom[3721] = 'b101001111;assign rom[3722] = 'b000111010;assign rom[3723] = 'b101110110;assign rom[3724] = 'b101100010;assign rom[3725] = 'b101001100;assign rom[3726] = 'b001001010;assign rom[3727] = 'b111011010;assign rom[3728] = 'b111011010;assign rom[3729] = 'b111011010;assign rom[3730] = 'b111011010;assign rom[3731] = 'b111011000;assign rom[3732] = 'b111011000;assign rom[3733] = 'b111011000;assign rom[3734] = 'b111011000;assign rom[3735] = 'b101111000;assign rom[3736] = 'b000110011;assign rom[3737] = 'b110000010;assign rom[3738] = 'b001101010;assign rom[3739] = 'b001011000;assign rom[3740] = 'b101001000;assign rom[3741] = 'b000101011;assign rom[3742] = 'b110000010;assign rom[3743] = 'b111000000;assign rom[3744] = 'b101001100;assign rom[3745] = 'b001001010;assign rom[3746] = 'b111111000;assign rom[3747] = 'b111101000;assign rom[3748] = 'b101001111;assign rom[3749] = 'b000111010;assign rom[3750] = 'b101110110;assign rom[3751] = 'b101100010;assign rom[3752] = 'b101001100;assign rom[3753] = 'b001001010;assign rom[3754] = 'b111011010;assign rom[3755] = 'b111011010;assign rom[3756] = 'b111011010;assign rom[3757] = 'b111011010;assign rom[3758] = 'b111011000;assign rom[3759] = 'b111011000;assign rom[3760] = 'b111011000;assign rom[3761] = 'b111011000;assign rom[3762] = 'b101111000;assign rom[3763] = 'b000110011;assign rom[3764] = 'b110000010;assign rom[3765] = 'b001101010;assign rom[3766] = 'b001011000;assign rom[3767] = 'b101001000;assign rom[3768] = 'b000101011;assign rom[3769] = 'b110000010;assign rom[3770] = 'b111000000;assign rom[3771] = 'b101001100;assign rom[3772] = 'b001001010;assign rom[3773] = 'b111111000;assign rom[3774] = 'b111101000;assign rom[3775] = 'b101001111;assign rom[3776] = 'b000111010;assign rom[3777] = 'b101110110;assign rom[3778] = 'b101100010;assign rom[3779] = 'b101001100;assign rom[3780] = 'b001001010;assign rom[3781] = 'b111011010;assign rom[3782] = 'b111011010;assign rom[3783] = 'b111011010;assign rom[3784] = 'b111011010;assign rom[3785] = 'b111011000;assign rom[3786] = 'b111011000;assign rom[3787] = 'b111011000;assign rom[3788] = 'b111011000;assign rom[3789] = 'b101111000;assign rom[3790] = 'b000110011;assign rom[3791] = 'b110000010;assign rom[3792] = 'b001101010;assign rom[3793] = 'b001011000;assign rom[3794] = 'b101001000;assign rom[3795] = 'b000101011;assign rom[3796] = 'b110000010;assign rom[3797] = 'b111000000;assign rom[3798] = 'b101001100;assign rom[3799] = 'b001001010;assign rom[3800] = 'b111111000;assign rom[3801] = 'b111101000;assign rom[3802] = 'b101001111;assign rom[3803] = 'b000111010;assign rom[3804] = 'b101110110;assign rom[3805] = 'b101100010;assign rom[3806] = 'b101001100;assign rom[3807] = 'b001001010;assign rom[3808] = 'b111011010;assign rom[3809] = 'b111011010;assign rom[3810] = 'b111011010;assign rom[3811] = 'b111011010;assign rom[3812] = 'b111011000;assign rom[3813] = 'b111011000;assign rom[3814] = 'b111011000;assign rom[3815] = 'b111011000;assign rom[3816] = 'b101111000;assign rom[3817] = 'b000110011;assign rom[3818] = 'b110000010;assign rom[3819] = 'b001101010;assign rom[3820] = 'b001011000;assign rom[3821] = 'b101001000;assign rom[3822] = 'b000101011;assign rom[3823] = 'b110000010;assign rom[3824] = 'b111000000;assign rom[3825] = 'b101001100;assign rom[3826] = 'b001001010;assign rom[3827] = 'b111111000;assign rom[3828] = 'b111101000;assign rom[3829] = 'b101001111;assign rom[3830] = 'b000111010;assign rom[3831] = 'b101110110;assign rom[3832] = 'b101100010;assign rom[3833] = 'b101001100;assign rom[3834] = 'b001001010;assign rom[3835] = 'b111011010;assign rom[3836] = 'b111011010;assign rom[3837] = 'b111011010;assign rom[3838] = 'b111011010;assign rom[3839] = 'b111011000;assign rom[3840] = 'b111011000;assign rom[3841] = 'b111011000;assign rom[3842] = 'b111011000;assign rom[3843] = 'b101111000;assign rom[3844] = 'b000110011;assign rom[3845] = 'b110000010;assign rom[3846] = 'b001101010;assign rom[3847] = 'b001011000;assign rom[3848] = 'b101001000;assign rom[3849] = 'b000101011;assign rom[3850] = 'b110000010;assign rom[3851] = 'b111000000;assign rom[3852] = 'b101001100;assign rom[3853] = 'b001001010;assign rom[3854] = 'b111111000;assign rom[3855] = 'b111101000;assign rom[3856] = 'b101001111;assign rom[3857] = 'b000111010;assign rom[3858] = 'b101110110;assign rom[3859] = 'b101100010;assign rom[3860] = 'b101001100;assign rom[3861] = 'b001001010;assign rom[3862] = 'b111011010;assign rom[3863] = 'b111011010;assign rom[3864] = 'b111011010;assign rom[3865] = 'b111011010;assign rom[3866] = 'b111011000;assign rom[3867] = 'b111011000;assign rom[3868] = 'b111011000;assign rom[3869] = 'b111011000;assign rom[3870] = 'b101111000;assign rom[3871] = 'b000110011;assign rom[3872] = 'b110000010;assign rom[3873] = 'b001101010;assign rom[3874] = 'b001011000;assign rom[3875] = 'b101001000;assign rom[3876] = 'b000101011;assign rom[3877] = 'b110000010;assign rom[3878] = 'b111000000;assign rom[3879] = 'b101001100;assign rom[3880] = 'b001001010;assign rom[3881] = 'b001000110;assign rom[3882] = 'b001100100;assign rom[3883] = 'b101100010;assign rom[3884] = 'b101001100;assign rom[3885] = 'b001001010;assign rom[3886] = 'b111011010;assign rom[3887] = 'b111011010;assign rom[3888] = 'b111011010;assign rom[3889] = 'b111011010;assign rom[3890] = 'b111011000;assign rom[3891] = 'b111011000;assign rom[3892] = 'b111011000;assign rom[3893] = 'b111011000;assign rom[3894] = 'b101111000;assign rom[3895] = 'b000110011;assign rom[3896] = 'b110000010;assign rom[3897] = 'b001101010;assign rom[3898] = 'b001011000;assign rom[3899] = 'b101001000;assign rom[3900] = 'b000101011;assign rom[3901] = 'b110000010;assign rom[3902] = 'b111000000;assign rom[3903] = 'b101001100;assign rom[3904] = 'b001001010;assign rom[3905] = 'b111111000;assign rom[3906] = 'b111101000;assign rom[3907] = 'b101001111;assign rom[3908] = 'b000111010;assign rom[3909] = 'b101110110;assign rom[3910] = 'b101100010;assign rom[3911] = 'b101001100;assign rom[3912] = 'b001001010;assign rom[3913] = 'b111011010;assign rom[3914] = 'b111011010;assign rom[3915] = 'b111011010;assign rom[3916] = 'b111011010;assign rom[3917] = 'b111011000;assign rom[3918] = 'b111011000;assign rom[3919] = 'b111011000;assign rom[3920] = 'b111011000;assign rom[3921] = 'b101111000;assign rom[3922] = 'b000110011;assign rom[3923] = 'b110000010;assign rom[3924] = 'b001101010;assign rom[3925] = 'b001011000;assign rom[3926] = 'b101001000;assign rom[3927] = 'b000101011;assign rom[3928] = 'b110000010;assign rom[3929] = 'b111000000;assign rom[3930] = 'b101001100;assign rom[3931] = 'b001001010;assign rom[3932] = 'b111111000;assign rom[3933] = 'b111101000;assign rom[3934] = 'b101001111;assign rom[3935] = 'b000111010;assign rom[3936] = 'b101110110;assign rom[3937] = 'b101100010;assign rom[3938] = 'b101001100;assign rom[3939] = 'b001001010;assign rom[3940] = 'b111011010;assign rom[3941] = 'b111011010;assign rom[3942] = 'b111011010;assign rom[3943] = 'b111011010;assign rom[3944] = 'b111011000;assign rom[3945] = 'b111011000;assign rom[3946] = 'b111011000;assign rom[3947] = 'b111011000;assign rom[3948] = 'b101111000;assign rom[3949] = 'b000110011;assign rom[3950] = 'b110000010;assign rom[3951] = 'b001101010;assign rom[3952] = 'b001011000;assign rom[3953] = 'b101001000;assign rom[3954] = 'b000101011;assign rom[3955] = 'b110000010;assign rom[3956] = 'b111000000;assign rom[3957] = 'b101001100;assign rom[3958] = 'b001001010;assign rom[3959] = 'b111111000;assign rom[3960] = 'b111101000;assign rom[3961] = 'b101001111;assign rom[3962] = 'b000111010;assign rom[3963] = 'b101110110;assign rom[3964] = 'b101100010;assign rom[3965] = 'b101001100;assign rom[3966] = 'b001001010;assign rom[3967] = 'b111011010;assign rom[3968] = 'b111011010;assign rom[3969] = 'b111011010;assign rom[3970] = 'b111011010;assign rom[3971] = 'b111011000;assign rom[3972] = 'b111011000;assign rom[3973] = 'b111011000;assign rom[3974] = 'b111011000;assign rom[3975] = 'b101111000;assign rom[3976] = 'b000110011;assign rom[3977] = 'b110000010;assign rom[3978] = 'b001101010;assign rom[3979] = 'b001011000;assign rom[3980] = 'b101001000;assign rom[3981] = 'b000101011;assign rom[3982] = 'b110000010;assign rom[3983] = 'b111000000;assign rom[3984] = 'b101001100;assign rom[3985] = 'b001001010;assign rom[3986] = 'b111111000;assign rom[3987] = 'b111101000;assign rom[3988] = 'b101001111;assign rom[3989] = 'b000111010;assign rom[3990] = 'b101110110;assign rom[3991] = 'b101100010;assign rom[3992] = 'b101001100;assign rom[3993] = 'b001001010;assign rom[3994] = 'b111011010;assign rom[3995] = 'b111011010;assign rom[3996] = 'b111011010;assign rom[3997] = 'b111011010;assign rom[3998] = 'b111011000;assign rom[3999] = 'b111011000;assign rom[4000] = 'b111011000;assign rom[4001] = 'b111011000;assign rom[4002] = 'b101111000;assign rom[4003] = 'b000110011;assign rom[4004] = 'b110000010;assign rom[4005] = 'b001101010;assign rom[4006] = 'b001011000;assign rom[4007] = 'b101001000;assign rom[4008] = 'b000101011;assign rom[4009] = 'b110000010;assign rom[4010] = 'b111000000;assign rom[4011] = 'b101001100;assign rom[4012] = 'b001001010;assign rom[4013] = 'b111111000;assign rom[4014] = 'b111101000;assign rom[4015] = 'b101001111;assign rom[4016] = 'b000111010;assign rom[4017] = 'b101110110;assign rom[4018] = 'b101100010;assign rom[4019] = 'b101001100;assign rom[4020] = 'b001001010;assign rom[4021] = 'b111011010;assign rom[4022] = 'b111011010;assign rom[4023] = 'b111011010;assign rom[4024] = 'b111011010;assign rom[4025] = 'b111011000;assign rom[4026] = 'b111011000;assign rom[4027] = 'b111011000;assign rom[4028] = 'b111011000;assign rom[4029] = 'b101111000;assign rom[4030] = 'b000110011;assign rom[4031] = 'b110000010;assign rom[4032] = 'b001101010;assign rom[4033] = 'b001011000;assign rom[4034] = 'b101001000;assign rom[4035] = 'b000101011;assign rom[4036] = 'b110000010;assign rom[4037] = 'b111000000;assign rom[4038] = 'b101001100;assign rom[4039] = 'b001001010;assign rom[4040] = 'b111111000;assign rom[4041] = 'b111101000;assign rom[4042] = 'b101001111;assign rom[4043] = 'b000111010;assign rom[4044] = 'b101110110;assign rom[4045] = 'b101100010;assign rom[4046] = 'b101001100;assign rom[4047] = 'b001001010;assign rom[4048] = 'b111011010;assign rom[4049] = 'b111011010;assign rom[4050] = 'b111011010;assign rom[4051] = 'b111011010;assign rom[4052] = 'b111011000;assign rom[4053] = 'b111011000;assign rom[4054] = 'b111011000;assign rom[4055] = 'b111011000;assign rom[4056] = 'b101111000;assign rom[4057] = 'b000110011;assign rom[4058] = 'b110000010;assign rom[4059] = 'b001101010;assign rom[4060] = 'b001011000;assign rom[4061] = 'b101001000;assign rom[4062] = 'b000101011;assign rom[4063] = 'b110000010;assign rom[4064] = 'b111000000;assign rom[4065] = 'b101001100;assign rom[4066] = 'b001001010;assign rom[4067] = 'b111111000;assign rom[4068] = 'b111101000;assign rom[4069] = 'b101001111;assign rom[4070] = 'b000111010;assign rom[4071] = 'b101110110;assign rom[4072] = 'b101100010;assign rom[4073] = 'b101001100;assign rom[4074] = 'b001001010;assign rom[4075] = 'b111011010;assign rom[4076] = 'b111011010;assign rom[4077] = 'b111011010;assign rom[4078] = 'b111011010;assign rom[4079] = 'b111011000;assign rom[4080] = 'b111011000;assign rom[4081] = 'b111011000;assign rom[4082] = 'b111011000;assign rom[4083] = 'b101111000;assign rom[4084] = 'b000110011;assign rom[4085] = 'b110000010;assign rom[4086] = 'b001101010;assign rom[4087] = 'b001011000;assign rom[4088] = 'b101001000;assign rom[4089] = 'b000101011;assign rom[4090] = 'b110000010;assign rom[4091] = 'b111000000;assign rom[4092] = 'b101001100;assign rom[4093] = 'b001001010;assign rom[4094] = 'b111111000;assign rom[4095] = 'b111101000;assign rom[4096] = 'b101001111;assign rom[4097] = 'b000111010;assign rom[4098] = 'b101110110;assign rom[4099] = 'b101100010;assign rom[4100] = 'b101001100;assign rom[4101] = 'b001001010;assign rom[4102] = 'b111011010;assign rom[4103] = 'b111011010;assign rom[4104] = 'b111011010;assign rom[4105] = 'b111011010;assign rom[4106] = 'b111011000;assign rom[4107] = 'b111011000;assign rom[4108] = 'b111011000;assign rom[4109] = 'b111011000;assign rom[4110] = 'b101111000;assign rom[4111] = 'b000110011;assign rom[4112] = 'b110000010;assign rom[4113] = 'b001101010;assign rom[4114] = 'b001011000;assign rom[4115] = 'b101001000;assign rom[4116] = 'b000101011;assign rom[4117] = 'b110000010;assign rom[4118] = 'b111000000;assign rom[4119] = 'b101001100;assign rom[4120] = 'b001001010;assign rom[4121] = 'b001000110;assign rom[4122] = 'b001100100;assign rom[4123] = 'b101100010;assign rom[4124] = 'b101001100;assign rom[4125] = 'b001001010;assign rom[4126] = 'b111011010;assign rom[4127] = 'b111011010;assign rom[4128] = 'b111011010;assign rom[4129] = 'b111011010;assign rom[4130] = 'b111011000;assign rom[4131] = 'b111011000;assign rom[4132] = 'b111011000;assign rom[4133] = 'b111011000;assign rom[4134] = 'b101111000;assign rom[4135] = 'b000110011;assign rom[4136] = 'b110000010;assign rom[4137] = 'b001101010;assign rom[4138] = 'b001011000;assign rom[4139] = 'b101001000;assign rom[4140] = 'b000101011;assign rom[4141] = 'b110000010;assign rom[4142] = 'b111000000;assign rom[4143] = 'b101001100;assign rom[4144] = 'b001001010;assign rom[4145] = 'b111111000;assign rom[4146] = 'b111101000;assign rom[4147] = 'b101001111;assign rom[4148] = 'b000111010;assign rom[4149] = 'b101110110;assign rom[4150] = 'b101100010;assign rom[4151] = 'b101001100;assign rom[4152] = 'b001001010;assign rom[4153] = 'b111011010;assign rom[4154] = 'b111011010;assign rom[4155] = 'b111011010;assign rom[4156] = 'b111011010;assign rom[4157] = 'b111011000;assign rom[4158] = 'b111011000;assign rom[4159] = 'b111011000;assign rom[4160] = 'b111011000;assign rom[4161] = 'b101111000;assign rom[4162] = 'b000110011;assign rom[4163] = 'b110000010;assign rom[4164] = 'b001101010;assign rom[4165] = 'b001011000;assign rom[4166] = 'b101001000;assign rom[4167] = 'b000101011;assign rom[4168] = 'b110000010;assign rom[4169] = 'b111000000;assign rom[4170] = 'b101001100;assign rom[4171] = 'b001001010;assign rom[4172] = 'b111111000;assign rom[4173] = 'b111101000;assign rom[4174] = 'b101001111;assign rom[4175] = 'b000111010;assign rom[4176] = 'b101110110;assign rom[4177] = 'b101100010;assign rom[4178] = 'b101001100;assign rom[4179] = 'b001001010;assign rom[4180] = 'b111011010;assign rom[4181] = 'b111011010;assign rom[4182] = 'b111011010;assign rom[4183] = 'b111011010;assign rom[4184] = 'b111011000;assign rom[4185] = 'b111011000;assign rom[4186] = 'b111011000;assign rom[4187] = 'b111011000;assign rom[4188] = 'b101111000;assign rom[4189] = 'b000110011;assign rom[4190] = 'b110000010;assign rom[4191] = 'b001101010;assign rom[4192] = 'b001011000;assign rom[4193] = 'b101001000;assign rom[4194] = 'b000101011;assign rom[4195] = 'b110000010;assign rom[4196] = 'b111000000;assign rom[4197] = 'b101001100;assign rom[4198] = 'b001001010;assign rom[4199] = 'b111111000;assign rom[4200] = 'b111101000;assign rom[4201] = 'b101001111;assign rom[4202] = 'b000111010;assign rom[4203] = 'b101110110;assign rom[4204] = 'b101100010;assign rom[4205] = 'b101001100;assign rom[4206] = 'b001001010;assign rom[4207] = 'b111011010;assign rom[4208] = 'b111011010;assign rom[4209] = 'b111011010;assign rom[4210] = 'b111011010;assign rom[4211] = 'b111011000;assign rom[4212] = 'b111011000;assign rom[4213] = 'b111011000;assign rom[4214] = 'b111011000;assign rom[4215] = 'b101111000;assign rom[4216] = 'b000110011;assign rom[4217] = 'b110000010;assign rom[4218] = 'b001101010;assign rom[4219] = 'b001011000;assign rom[4220] = 'b101001000;assign rom[4221] = 'b000101011;assign rom[4222] = 'b110000010;assign rom[4223] = 'b111000000;assign rom[4224] = 'b101001100;assign rom[4225] = 'b001001010;assign rom[4226] = 'b111111000;assign rom[4227] = 'b111101000;assign rom[4228] = 'b101001111;assign rom[4229] = 'b000111010;assign rom[4230] = 'b101110110;assign rom[4231] = 'b101100010;assign rom[4232] = 'b101001100;assign rom[4233] = 'b001001010;assign rom[4234] = 'b111011010;assign rom[4235] = 'b111011010;assign rom[4236] = 'b111011010;assign rom[4237] = 'b111011010;assign rom[4238] = 'b111011000;assign rom[4239] = 'b111011000;assign rom[4240] = 'b111011000;assign rom[4241] = 'b111011000;assign rom[4242] = 'b101111000;assign rom[4243] = 'b000110011;assign rom[4244] = 'b110000010;assign rom[4245] = 'b001101010;assign rom[4246] = 'b001011000;assign rom[4247] = 'b101001000;assign rom[4248] = 'b000101011;assign rom[4249] = 'b110000010;assign rom[4250] = 'b111000000;assign rom[4251] = 'b101001100;assign rom[4252] = 'b001001010;assign rom[4253] = 'b111111000;assign rom[4254] = 'b111101000;assign rom[4255] = 'b101001111;assign rom[4256] = 'b000111010;assign rom[4257] = 'b101110110;assign rom[4258] = 'b101100010;assign rom[4259] = 'b101001100;assign rom[4260] = 'b001001010;assign rom[4261] = 'b111011010;assign rom[4262] = 'b111011010;assign rom[4263] = 'b111011010;assign rom[4264] = 'b111011010;assign rom[4265] = 'b111011000;assign rom[4266] = 'b111011000;assign rom[4267] = 'b111011000;assign rom[4268] = 'b111011000;assign rom[4269] = 'b101111000;assign rom[4270] = 'b000110011;assign rom[4271] = 'b110000010;assign rom[4272] = 'b001101010;assign rom[4273] = 'b001011000;assign rom[4274] = 'b101001000;assign rom[4275] = 'b000101011;assign rom[4276] = 'b110000010;assign rom[4277] = 'b111000000;assign rom[4278] = 'b101001100;assign rom[4279] = 'b001001010;assign rom[4280] = 'b111111000;assign rom[4281] = 'b111101000;assign rom[4282] = 'b101001111;assign rom[4283] = 'b000111010;assign rom[4284] = 'b101110110;assign rom[4285] = 'b101100010;assign rom[4286] = 'b101001100;assign rom[4287] = 'b001001010;assign rom[4288] = 'b111011010;assign rom[4289] = 'b111011010;assign rom[4290] = 'b111011010;assign rom[4291] = 'b111011010;assign rom[4292] = 'b111011000;assign rom[4293] = 'b111011000;assign rom[4294] = 'b111011000;assign rom[4295] = 'b111011000;assign rom[4296] = 'b101111000;assign rom[4297] = 'b000110011;assign rom[4298] = 'b110000010;assign rom[4299] = 'b001101010;assign rom[4300] = 'b001011000;assign rom[4301] = 'b101001000;assign rom[4302] = 'b000101011;assign rom[4303] = 'b110000010;assign rom[4304] = 'b111000000;assign rom[4305] = 'b101001100;assign rom[4306] = 'b001001010;assign rom[4307] = 'b111111000;assign rom[4308] = 'b111101000;assign rom[4309] = 'b101001111;assign rom[4310] = 'b000111010;assign rom[4311] = 'b101110110;assign rom[4312] = 'b101100010;assign rom[4313] = 'b101001100;assign rom[4314] = 'b001001010;assign rom[4315] = 'b111011010;assign rom[4316] = 'b111011010;assign rom[4317] = 'b111011010;assign rom[4318] = 'b111011010;assign rom[4319] = 'b111011000;assign rom[4320] = 'b111011000;assign rom[4321] = 'b111011000;assign rom[4322] = 'b111011000;assign rom[4323] = 'b101111000;assign rom[4324] = 'b000110011;assign rom[4325] = 'b110000010;assign rom[4326] = 'b001101010;assign rom[4327] = 'b001011000;assign rom[4328] = 'b101001000;assign rom[4329] = 'b000101011;assign rom[4330] = 'b110000010;assign rom[4331] = 'b111000000;assign rom[4332] = 'b101001100;assign rom[4333] = 'b001001010;assign rom[4334] = 'b111111000;assign rom[4335] = 'b111101000;assign rom[4336] = 'b101001111;assign rom[4337] = 'b000111010;assign rom[4338] = 'b101110110;assign rom[4339] = 'b101100010;assign rom[4340] = 'b101001100;assign rom[4341] = 'b001001010;assign rom[4342] = 'b111011010;assign rom[4343] = 'b111011010;assign rom[4344] = 'b111011010;assign rom[4345] = 'b111011010;assign rom[4346] = 'b111011000;assign rom[4347] = 'b111011000;assign rom[4348] = 'b111011000;assign rom[4349] = 'b111011000;assign rom[4350] = 'b101111000;assign rom[4351] = 'b000110011;assign rom[4352] = 'b110000010;assign rom[4353] = 'b001101010;assign rom[4354] = 'b001011000;assign rom[4355] = 'b101001000;assign rom[4356] = 'b000101011;assign rom[4357] = 'b110000010;assign rom[4358] = 'b111000000;assign rom[4359] = 'b101001100;assign rom[4360] = 'b001001010;assign rom[4361] = 'b001000110;assign rom[4362] = 'b001100100;assign rom[4363] = 'b101100010;assign rom[4364] = 'b101001100;assign rom[4365] = 'b001001010;assign rom[4366] = 'b111011010;assign rom[4367] = 'b111011010;assign rom[4368] = 'b111011010;assign rom[4369] = 'b111011010;assign rom[4370] = 'b111011000;assign rom[4371] = 'b111011000;assign rom[4372] = 'b111011000;assign rom[4373] = 'b111011000;assign rom[4374] = 'b101111000;assign rom[4375] = 'b000110011;assign rom[4376] = 'b110000010;assign rom[4377] = 'b001101010;assign rom[4378] = 'b001011000;assign rom[4379] = 'b101001000;assign rom[4380] = 'b000101011;assign rom[4381] = 'b110000010;assign rom[4382] = 'b111000000;assign rom[4383] = 'b101001100;assign rom[4384] = 'b001001010;assign rom[4385] = 'b111111000;assign rom[4386] = 'b111101000;assign rom[4387] = 'b101001111;assign rom[4388] = 'b000111010;assign rom[4389] = 'b101110110;assign rom[4390] = 'b101100010;assign rom[4391] = 'b101001100;assign rom[4392] = 'b001001010;assign rom[4393] = 'b111011010;assign rom[4394] = 'b111011010;assign rom[4395] = 'b111011010;assign rom[4396] = 'b111011010;assign rom[4397] = 'b111011000;assign rom[4398] = 'b111011000;assign rom[4399] = 'b111011000;assign rom[4400] = 'b111011000;assign rom[4401] = 'b101111000;assign rom[4402] = 'b000110011;assign rom[4403] = 'b110000010;assign rom[4404] = 'b001101010;assign rom[4405] = 'b001011000;assign rom[4406] = 'b101001000;assign rom[4407] = 'b000101011;assign rom[4408] = 'b110000010;assign rom[4409] = 'b111000000;assign rom[4410] = 'b101001100;assign rom[4411] = 'b001001010;assign rom[4412] = 'b111111000;assign rom[4413] = 'b111101000;assign rom[4414] = 'b101001111;assign rom[4415] = 'b000111010;assign rom[4416] = 'b101110110;assign rom[4417] = 'b101100010;assign rom[4418] = 'b101001100;assign rom[4419] = 'b001001010;assign rom[4420] = 'b111011010;assign rom[4421] = 'b111011010;assign rom[4422] = 'b111011010;assign rom[4423] = 'b111011010;assign rom[4424] = 'b111011000;assign rom[4425] = 'b111011000;assign rom[4426] = 'b111011000;assign rom[4427] = 'b111011000;assign rom[4428] = 'b101111000;assign rom[4429] = 'b000110011;assign rom[4430] = 'b110000010;assign rom[4431] = 'b001101010;assign rom[4432] = 'b001011000;assign rom[4433] = 'b101001000;assign rom[4434] = 'b000101011;assign rom[4435] = 'b110000010;assign rom[4436] = 'b111000000;assign rom[4437] = 'b101001100;assign rom[4438] = 'b001001010;assign rom[4439] = 'b111111000;assign rom[4440] = 'b111101000;assign rom[4441] = 'b101001111;assign rom[4442] = 'b000111010;assign rom[4443] = 'b101110110;assign rom[4444] = 'b101100010;assign rom[4445] = 'b101001100;assign rom[4446] = 'b001001010;assign rom[4447] = 'b111011010;assign rom[4448] = 'b111011010;assign rom[4449] = 'b111011010;assign rom[4450] = 'b111011010;assign rom[4451] = 'b111011000;assign rom[4452] = 'b111011000;assign rom[4453] = 'b111011000;assign rom[4454] = 'b111011000;assign rom[4455] = 'b101111000;assign rom[4456] = 'b000110011;assign rom[4457] = 'b110000010;assign rom[4458] = 'b001101010;assign rom[4459] = 'b001011000;assign rom[4460] = 'b101001000;assign rom[4461] = 'b000101011;assign rom[4462] = 'b110000010;assign rom[4463] = 'b111000000;assign rom[4464] = 'b101001100;assign rom[4465] = 'b001001010;assign rom[4466] = 'b111111000;assign rom[4467] = 'b111101000;assign rom[4468] = 'b101001111;assign rom[4469] = 'b000111010;assign rom[4470] = 'b101110110;assign rom[4471] = 'b101100010;assign rom[4472] = 'b101001100;assign rom[4473] = 'b001001010;assign rom[4474] = 'b111011010;assign rom[4475] = 'b111011010;assign rom[4476] = 'b111011010;assign rom[4477] = 'b111011010;assign rom[4478] = 'b111011000;assign rom[4479] = 'b111011000;assign rom[4480] = 'b111011000;assign rom[4481] = 'b111011000;assign rom[4482] = 'b101111000;assign rom[4483] = 'b000110011;assign rom[4484] = 'b110000010;assign rom[4485] = 'b001101010;assign rom[4486] = 'b001011000;assign rom[4487] = 'b101001000;assign rom[4488] = 'b000101011;assign rom[4489] = 'b110000010;assign rom[4490] = 'b111000000;assign rom[4491] = 'b101001100;assign rom[4492] = 'b001001010;assign rom[4493] = 'b111111000;assign rom[4494] = 'b111101000;assign rom[4495] = 'b101001111;assign rom[4496] = 'b000111010;assign rom[4497] = 'b101110110;assign rom[4498] = 'b101100010;assign rom[4499] = 'b101001100;assign rom[4500] = 'b001001010;assign rom[4501] = 'b111011010;assign rom[4502] = 'b111011010;assign rom[4503] = 'b111011010;assign rom[4504] = 'b111011010;assign rom[4505] = 'b111011000;assign rom[4506] = 'b111011000;assign rom[4507] = 'b111011000;assign rom[4508] = 'b111011000;assign rom[4509] = 'b101111000;assign rom[4510] = 'b000110011;assign rom[4511] = 'b110000010;assign rom[4512] = 'b001101010;assign rom[4513] = 'b001011000;assign rom[4514] = 'b101001000;assign rom[4515] = 'b000101011;assign rom[4516] = 'b110000010;assign rom[4517] = 'b111000000;assign rom[4518] = 'b101001100;assign rom[4519] = 'b001001010;assign rom[4520] = 'b111111000;assign rom[4521] = 'b111101000;assign rom[4522] = 'b101001111;assign rom[4523] = 'b000111010;assign rom[4524] = 'b101110110;assign rom[4525] = 'b101100010;assign rom[4526] = 'b101001100;assign rom[4527] = 'b001001010;assign rom[4528] = 'b111011010;assign rom[4529] = 'b111011010;assign rom[4530] = 'b111011010;assign rom[4531] = 'b111011010;assign rom[4532] = 'b111011000;assign rom[4533] = 'b111011000;assign rom[4534] = 'b111011000;assign rom[4535] = 'b111011000;assign rom[4536] = 'b101111000;assign rom[4537] = 'b000110011;assign rom[4538] = 'b110000010;assign rom[4539] = 'b001101010;assign rom[4540] = 'b001011000;assign rom[4541] = 'b101001000;assign rom[4542] = 'b000101011;assign rom[4543] = 'b110000010;assign rom[4544] = 'b111000000;assign rom[4545] = 'b101001100;assign rom[4546] = 'b001001010;assign rom[4547] = 'b111111000;assign rom[4548] = 'b111101000;assign rom[4549] = 'b101001111;assign rom[4550] = 'b000111010;assign rom[4551] = 'b101110110;assign rom[4552] = 'b101100010;assign rom[4553] = 'b101001100;assign rom[4554] = 'b001001010;assign rom[4555] = 'b111011010;assign rom[4556] = 'b111011010;assign rom[4557] = 'b111011010;assign rom[4558] = 'b111011010;assign rom[4559] = 'b111011000;assign rom[4560] = 'b111011000;assign rom[4561] = 'b111011000;assign rom[4562] = 'b111011000;assign rom[4563] = 'b101111000;assign rom[4564] = 'b000110011;assign rom[4565] = 'b110000010;assign rom[4566] = 'b001101010;assign rom[4567] = 'b001011000;assign rom[4568] = 'b101001000;assign rom[4569] = 'b000101011;assign rom[4570] = 'b110000010;assign rom[4571] = 'b111000000;assign rom[4572] = 'b101001100;assign rom[4573] = 'b001001010;assign rom[4574] = 'b111111000;assign rom[4575] = 'b111101000;assign rom[4576] = 'b101001111;assign rom[4577] = 'b000111010;assign rom[4578] = 'b101110110;assign rom[4579] = 'b101100010;assign rom[4580] = 'b101001100;assign rom[4581] = 'b001001010;assign rom[4582] = 'b111011010;assign rom[4583] = 'b111011010;assign rom[4584] = 'b111011010;assign rom[4585] = 'b111011010;assign rom[4586] = 'b111011000;assign rom[4587] = 'b111011000;assign rom[4588] = 'b111011000;assign rom[4589] = 'b111011000;assign rom[4590] = 'b101111000;assign rom[4591] = 'b000110011;assign rom[4592] = 'b110000010;assign rom[4593] = 'b001101010;assign rom[4594] = 'b001011000;assign rom[4595] = 'b101001000;assign rom[4596] = 'b000101011;assign rom[4597] = 'b110000010;assign rom[4598] = 'b111000000;assign rom[4599] = 'b101001100;assign rom[4600] = 'b001001010;assign rom[4601] = 'b001000110;assign rom[4602] = 'b001100100;assign rom[4603] = 'b101100010;assign rom[4604] = 'b101001100;assign rom[4605] = 'b001001010;assign rom[4606] = 'b111011010;assign rom[4607] = 'b111011010;assign rom[4608] = 'b111011010;assign rom[4609] = 'b111011010;assign rom[4610] = 'b111011000;assign rom[4611] = 'b111011000;assign rom[4612] = 'b111011000;assign rom[4613] = 'b111011000;assign rom[4614] = 'b101111000;assign rom[4615] = 'b000110011;assign rom[4616] = 'b110000010;assign rom[4617] = 'b001101010;assign rom[4618] = 'b001011000;assign rom[4619] = 'b101001000;assign rom[4620] = 'b000101011;assign rom[4621] = 'b110000010;assign rom[4622] = 'b111000000;assign rom[4623] = 'b101001100;assign rom[4624] = 'b001001010;assign rom[4625] = 'b111111000;assign rom[4626] = 'b111101000;assign rom[4627] = 'b101001111;assign rom[4628] = 'b000111010;assign rom[4629] = 'b101110110;assign rom[4630] = 'b101100010;assign rom[4631] = 'b101001100;assign rom[4632] = 'b001001010;assign rom[4633] = 'b111011010;assign rom[4634] = 'b111011010;assign rom[4635] = 'b111011010;assign rom[4636] = 'b111011010;assign rom[4637] = 'b111011000;assign rom[4638] = 'b111011000;assign rom[4639] = 'b111011000;assign rom[4640] = 'b111011000;assign rom[4641] = 'b101111000;assign rom[4642] = 'b000110011;assign rom[4643] = 'b110000010;assign rom[4644] = 'b001101010;assign rom[4645] = 'b001011000;assign rom[4646] = 'b101001000;assign rom[4647] = 'b000101011;assign rom[4648] = 'b110000010;assign rom[4649] = 'b111000000;assign rom[4650] = 'b101001100;assign rom[4651] = 'b001001010;assign rom[4652] = 'b111111000;assign rom[4653] = 'b111101000;assign rom[4654] = 'b101001111;assign rom[4655] = 'b000111010;assign rom[4656] = 'b101110110;assign rom[4657] = 'b101100010;assign rom[4658] = 'b101001100;assign rom[4659] = 'b001001010;assign rom[4660] = 'b111011010;assign rom[4661] = 'b111011010;assign rom[4662] = 'b111011010;assign rom[4663] = 'b111011010;assign rom[4664] = 'b111011000;assign rom[4665] = 'b111011000;assign rom[4666] = 'b111011000;assign rom[4667] = 'b111011000;assign rom[4668] = 'b101111000;assign rom[4669] = 'b000110011;assign rom[4670] = 'b110000010;assign rom[4671] = 'b001101010;assign rom[4672] = 'b001011000;assign rom[4673] = 'b101001000;assign rom[4674] = 'b000101011;assign rom[4675] = 'b110000010;assign rom[4676] = 'b111000000;assign rom[4677] = 'b101001100;assign rom[4678] = 'b001001010;assign rom[4679] = 'b111111000;assign rom[4680] = 'b111101000;assign rom[4681] = 'b101001111;assign rom[4682] = 'b000111010;assign rom[4683] = 'b101110110;assign rom[4684] = 'b101100010;assign rom[4685] = 'b101001100;assign rom[4686] = 'b001001010;assign rom[4687] = 'b111011010;assign rom[4688] = 'b111011010;assign rom[4689] = 'b111011010;assign rom[4690] = 'b111011010;assign rom[4691] = 'b111011000;assign rom[4692] = 'b111011000;assign rom[4693] = 'b111011000;assign rom[4694] = 'b111011000;assign rom[4695] = 'b101111000;assign rom[4696] = 'b000110011;assign rom[4697] = 'b110000010;assign rom[4698] = 'b001101010;assign rom[4699] = 'b001011000;assign rom[4700] = 'b101001000;assign rom[4701] = 'b000101011;assign rom[4702] = 'b110000010;assign rom[4703] = 'b111000000;assign rom[4704] = 'b101001100;assign rom[4705] = 'b001001010;assign rom[4706] = 'b111111000;assign rom[4707] = 'b111101000;assign rom[4708] = 'b101001111;assign rom[4709] = 'b000111010;assign rom[4710] = 'b101110110;assign rom[4711] = 'b101100010;assign rom[4712] = 'b101001100;assign rom[4713] = 'b001001010;assign rom[4714] = 'b111011010;assign rom[4715] = 'b111011010;assign rom[4716] = 'b111011010;assign rom[4717] = 'b111011010;assign rom[4718] = 'b111011000;assign rom[4719] = 'b111011000;assign rom[4720] = 'b111011000;assign rom[4721] = 'b111011000;assign rom[4722] = 'b101111000;assign rom[4723] = 'b000110011;assign rom[4724] = 'b110000010;assign rom[4725] = 'b001101010;assign rom[4726] = 'b001011000;assign rom[4727] = 'b101001000;assign rom[4728] = 'b000101011;assign rom[4729] = 'b110000010;assign rom[4730] = 'b111000000;assign rom[4731] = 'b101001100;assign rom[4732] = 'b001001010;assign rom[4733] = 'b111111000;assign rom[4734] = 'b111101000;assign rom[4735] = 'b101001111;assign rom[4736] = 'b000111010;assign rom[4737] = 'b101110110;assign rom[4738] = 'b101100010;assign rom[4739] = 'b101001100;assign rom[4740] = 'b001001010;assign rom[4741] = 'b111011010;assign rom[4742] = 'b111011010;assign rom[4743] = 'b111011010;assign rom[4744] = 'b111011010;assign rom[4745] = 'b111011000;assign rom[4746] = 'b111011000;assign rom[4747] = 'b111011000;assign rom[4748] = 'b111011000;assign rom[4749] = 'b101111000;assign rom[4750] = 'b000110011;assign rom[4751] = 'b110000010;assign rom[4752] = 'b001101010;assign rom[4753] = 'b001011000;assign rom[4754] = 'b101001000;assign rom[4755] = 'b000101011;assign rom[4756] = 'b110000010;assign rom[4757] = 'b111000000;assign rom[4758] = 'b101001100;assign rom[4759] = 'b001001010;assign rom[4760] = 'b111111000;assign rom[4761] = 'b111101000;assign rom[4762] = 'b101001111;assign rom[4763] = 'b000111010;assign rom[4764] = 'b101110110;assign rom[4765] = 'b101100010;assign rom[4766] = 'b101001100;assign rom[4767] = 'b001001010;assign rom[4768] = 'b111011010;assign rom[4769] = 'b111011010;assign rom[4770] = 'b111011010;assign rom[4771] = 'b111011010;assign rom[4772] = 'b111011000;assign rom[4773] = 'b111011000;assign rom[4774] = 'b111011000;assign rom[4775] = 'b111011000;assign rom[4776] = 'b101111000;assign rom[4777] = 'b000110011;assign rom[4778] = 'b110000010;assign rom[4779] = 'b001101010;assign rom[4780] = 'b001011000;assign rom[4781] = 'b101001000;assign rom[4782] = 'b000101011;assign rom[4783] = 'b110000010;assign rom[4784] = 'b111000000;assign rom[4785] = 'b101001100;assign rom[4786] = 'b001001010;assign rom[4787] = 'b111111000;assign rom[4788] = 'b111101000;assign rom[4789] = 'b101001111;assign rom[4790] = 'b000111010;assign rom[4791] = 'b101110110;assign rom[4792] = 'b101100010;assign rom[4793] = 'b101001100;assign rom[4794] = 'b001001010;assign rom[4795] = 'b111011010;assign rom[4796] = 'b111011010;assign rom[4797] = 'b111011010;assign rom[4798] = 'b111011010;assign rom[4799] = 'b111011000;assign rom[4800] = 'b111011000;assign rom[4801] = 'b111011000;assign rom[4802] = 'b111011000;assign rom[4803] = 'b101111000;assign rom[4804] = 'b000110011;assign rom[4805] = 'b110000010;assign rom[4806] = 'b001101010;assign rom[4807] = 'b001011000;assign rom[4808] = 'b101001000;assign rom[4809] = 'b000101011;assign rom[4810] = 'b110000010;assign rom[4811] = 'b111000000;assign rom[4812] = 'b101001100;assign rom[4813] = 'b001001010;assign rom[4814] = 'b111111000;assign rom[4815] = 'b111101000;assign rom[4816] = 'b101001111;assign rom[4817] = 'b000111010;assign rom[4818] = 'b101110110;assign rom[4819] = 'b101100010;assign rom[4820] = 'b101001100;assign rom[4821] = 'b001001010;assign rom[4822] = 'b111011010;assign rom[4823] = 'b111011010;assign rom[4824] = 'b111011010;assign rom[4825] = 'b111011010;assign rom[4826] = 'b111011000;assign rom[4827] = 'b111011000;assign rom[4828] = 'b111011000;assign rom[4829] = 'b111011000;assign rom[4830] = 'b101111000;assign rom[4831] = 'b000110011;assign rom[4832] = 'b110000010;assign rom[4833] = 'b001101010;assign rom[4834] = 'b001011000;assign rom[4835] = 'b101001000;assign rom[4836] = 'b000101011;assign rom[4837] = 'b110000010;assign rom[4838] = 'b111000000;assign rom[4839] = 'b101001100;assign rom[4840] = 'b001001010;assign rom[4841] = 'b001000110;assign rom[4842] = 'b001100100;assign rom[4843] = 'b101100010;assign rom[4844] = 'b101001100;assign rom[4845] = 'b001001010;assign rom[4846] = 'b111011010;assign rom[4847] = 'b111011010;assign rom[4848] = 'b111011010;assign rom[4849] = 'b111011010;assign rom[4850] = 'b111011000;assign rom[4851] = 'b111011000;assign rom[4852] = 'b111011000;assign rom[4853] = 'b111011000;assign rom[4854] = 'b101111000;assign rom[4855] = 'b000110011;assign rom[4856] = 'b110000010;assign rom[4857] = 'b001101010;assign rom[4858] = 'b001011000;assign rom[4859] = 'b101001000;assign rom[4860] = 'b000101011;assign rom[4861] = 'b110000010;assign rom[4862] = 'b111000000;assign rom[4863] = 'b101001100;assign rom[4864] = 'b001001010;assign rom[4865] = 'b111111000;assign rom[4866] = 'b111101000;assign rom[4867] = 'b101001111;assign rom[4868] = 'b000111010;assign rom[4869] = 'b101110110;assign rom[4870] = 'b101100010;assign rom[4871] = 'b101001100;assign rom[4872] = 'b001001010;assign rom[4873] = 'b111011010;assign rom[4874] = 'b111011010;assign rom[4875] = 'b111011010;assign rom[4876] = 'b111011010;assign rom[4877] = 'b111011000;assign rom[4878] = 'b111011000;assign rom[4879] = 'b111011000;assign rom[4880] = 'b111011000;assign rom[4881] = 'b101111000;assign rom[4882] = 'b000110011;assign rom[4883] = 'b110000010;assign rom[4884] = 'b001101010;assign rom[4885] = 'b001011000;assign rom[4886] = 'b101001000;assign rom[4887] = 'b000101011;assign rom[4888] = 'b110000010;assign rom[4889] = 'b111000000;assign rom[4890] = 'b101001100;assign rom[4891] = 'b001001010;assign rom[4892] = 'b111111000;assign rom[4893] = 'b111101000;assign rom[4894] = 'b101001111;assign rom[4895] = 'b000111010;assign rom[4896] = 'b101110110;assign rom[4897] = 'b101100010;assign rom[4898] = 'b101001100;assign rom[4899] = 'b001001010;assign rom[4900] = 'b111011010;assign rom[4901] = 'b111011010;assign rom[4902] = 'b111011010;assign rom[4903] = 'b111011010;assign rom[4904] = 'b111011000;assign rom[4905] = 'b111011000;assign rom[4906] = 'b111011000;assign rom[4907] = 'b111011000;assign rom[4908] = 'b101111000;assign rom[4909] = 'b000110011;assign rom[4910] = 'b110000010;assign rom[4911] = 'b001101010;assign rom[4912] = 'b001011000;assign rom[4913] = 'b101001000;assign rom[4914] = 'b000101011;assign rom[4915] = 'b110000010;assign rom[4916] = 'b111000000;assign rom[4917] = 'b101001100;assign rom[4918] = 'b001001010;assign rom[4919] = 'b111111000;assign rom[4920] = 'b111101000;assign rom[4921] = 'b101001111;assign rom[4922] = 'b000111010;assign rom[4923] = 'b101110110;assign rom[4924] = 'b101100010;assign rom[4925] = 'b101001100;assign rom[4926] = 'b001001010;assign rom[4927] = 'b111011010;assign rom[4928] = 'b111011010;assign rom[4929] = 'b111011010;assign rom[4930] = 'b111011010;assign rom[4931] = 'b111011000;assign rom[4932] = 'b111011000;assign rom[4933] = 'b111011000;assign rom[4934] = 'b111011000;assign rom[4935] = 'b101111000;assign rom[4936] = 'b000110011;assign rom[4937] = 'b110000010;assign rom[4938] = 'b001101010;assign rom[4939] = 'b001011000;assign rom[4940] = 'b101001000;assign rom[4941] = 'b000101011;assign rom[4942] = 'b110000010;assign rom[4943] = 'b111000000;assign rom[4944] = 'b101001100;assign rom[4945] = 'b001001010;assign rom[4946] = 'b111111000;assign rom[4947] = 'b111101000;assign rom[4948] = 'b101001111;assign rom[4949] = 'b000111010;assign rom[4950] = 'b101110110;assign rom[4951] = 'b101100010;assign rom[4952] = 'b101001100;assign rom[4953] = 'b001001010;assign rom[4954] = 'b111011010;assign rom[4955] = 'b111011010;assign rom[4956] = 'b111011010;assign rom[4957] = 'b111011010;assign rom[4958] = 'b111011000;assign rom[4959] = 'b111011000;assign rom[4960] = 'b111011000;assign rom[4961] = 'b111011000;assign rom[4962] = 'b101111000;assign rom[4963] = 'b000110011;assign rom[4964] = 'b110000010;assign rom[4965] = 'b001101010;assign rom[4966] = 'b001011000;assign rom[4967] = 'b101001000;assign rom[4968] = 'b000101011;assign rom[4969] = 'b110000010;assign rom[4970] = 'b111000000;assign rom[4971] = 'b101001100;assign rom[4972] = 'b001001010;assign rom[4973] = 'b111111000;assign rom[4974] = 'b111101000;assign rom[4975] = 'b101001111;assign rom[4976] = 'b000111010;assign rom[4977] = 'b101110110;assign rom[4978] = 'b101100010;assign rom[4979] = 'b101001100;assign rom[4980] = 'b001001010;assign rom[4981] = 'b111011010;assign rom[4982] = 'b111011010;assign rom[4983] = 'b111011010;assign rom[4984] = 'b111011010;assign rom[4985] = 'b111011000;assign rom[4986] = 'b111011000;assign rom[4987] = 'b111011000;assign rom[4988] = 'b111011000;assign rom[4989] = 'b101111000;assign rom[4990] = 'b000110011;assign rom[4991] = 'b110000010;assign rom[4992] = 'b001101010;assign rom[4993] = 'b001011000;assign rom[4994] = 'b101001000;assign rom[4995] = 'b000101011;assign rom[4996] = 'b110000010;assign rom[4997] = 'b111000000;assign rom[4998] = 'b101001100;assign rom[4999] = 'b001001010;assign rom[5000] = 'b111111000;assign rom[5001] = 'b111101000;assign rom[5002] = 'b101001111;assign rom[5003] = 'b000111010;assign rom[5004] = 'b101110110;assign rom[5005] = 'b101100010;assign rom[5006] = 'b101001100;assign rom[5007] = 'b001001010;assign rom[5008] = 'b111011010;assign rom[5009] = 'b111011010;assign rom[5010] = 'b111011010;assign rom[5011] = 'b111011010;assign rom[5012] = 'b111011000;assign rom[5013] = 'b111011000;assign rom[5014] = 'b111011000;assign rom[5015] = 'b111011000;assign rom[5016] = 'b101111000;assign rom[5017] = 'b000110011;assign rom[5018] = 'b110000010;assign rom[5019] = 'b001101010;assign rom[5020] = 'b001011000;assign rom[5021] = 'b101001000;assign rom[5022] = 'b000101011;assign rom[5023] = 'b110000010;assign rom[5024] = 'b111000000;assign rom[5025] = 'b101001100;assign rom[5026] = 'b001001010;assign rom[5027] = 'b111111000;assign rom[5028] = 'b111101000;assign rom[5029] = 'b101001111;assign rom[5030] = 'b000111010;assign rom[5031] = 'b101110110;assign rom[5032] = 'b101100010;assign rom[5033] = 'b101001100;assign rom[5034] = 'b001001010;assign rom[5035] = 'b111011010;assign rom[5036] = 'b111011010;assign rom[5037] = 'b111011010;assign rom[5038] = 'b111011010;assign rom[5039] = 'b111011000;assign rom[5040] = 'b111011000;assign rom[5041] = 'b111011000;assign rom[5042] = 'b111011000;assign rom[5043] = 'b101111000;assign rom[5044] = 'b000110011;assign rom[5045] = 'b110000010;assign rom[5046] = 'b001101010;assign rom[5047] = 'b001011000;assign rom[5048] = 'b101001000;assign rom[5049] = 'b000101011;assign rom[5050] = 'b110000010;assign rom[5051] = 'b111000000;assign rom[5052] = 'b101001100;assign rom[5053] = 'b001001010;assign rom[5054] = 'b111111000;assign rom[5055] = 'b111101000;assign rom[5056] = 'b101001111;assign rom[5057] = 'b000111010;assign rom[5058] = 'b101110110;assign rom[5059] = 'b101100010;assign rom[5060] = 'b101001100;assign rom[5061] = 'b001001010;assign rom[5062] = 'b111011010;assign rom[5063] = 'b111011010;assign rom[5064] = 'b111011010;assign rom[5065] = 'b111011010;assign rom[5066] = 'b111011000;assign rom[5067] = 'b111011000;assign rom[5068] = 'b111011000;assign rom[5069] = 'b111011000;assign rom[5070] = 'b101111000;assign rom[5071] = 'b000110011;assign rom[5072] = 'b110000010;assign rom[5073] = 'b001101010;assign rom[5074] = 'b001011000;assign rom[5075] = 'b101001000;assign rom[5076] = 'b000101011;assign rom[5077] = 'b110000010;assign rom[5078] = 'b111000000;assign rom[5079] = 'b101001100;assign rom[5080] = 'b001001010;assign rom[5081] = 'b001000110;assign rom[5082] = 'b001100100;assign rom[5083] = 'b101100010;assign rom[5084] = 'b101001100;assign rom[5085] = 'b001001010;assign rom[5086] = 'b111011010;assign rom[5087] = 'b111011010;assign rom[5088] = 'b111011010;assign rom[5089] = 'b111011010;assign rom[5090] = 'b111011000;assign rom[5091] = 'b111011000;assign rom[5092] = 'b111011000;assign rom[5093] = 'b111011000;assign rom[5094] = 'b101111000;assign rom[5095] = 'b000110011;assign rom[5096] = 'b110000010;assign rom[5097] = 'b001101010;assign rom[5098] = 'b001011000;assign rom[5099] = 'b101001000;assign rom[5100] = 'b000101011;assign rom[5101] = 'b110000010;assign rom[5102] = 'b111000000;assign rom[5103] = 'b101001100;assign rom[5104] = 'b001001010;assign rom[5105] = 'b111111000;assign rom[5106] = 'b111101000;assign rom[5107] = 'b101001111;assign rom[5108] = 'b000111010;assign rom[5109] = 'b101110110;assign rom[5110] = 'b101100010;assign rom[5111] = 'b101001100;assign rom[5112] = 'b001001010;assign rom[5113] = 'b111011010;assign rom[5114] = 'b111011010;assign rom[5115] = 'b111011010;assign rom[5116] = 'b111011010;assign rom[5117] = 'b111011000;assign rom[5118] = 'b111011000;assign rom[5119] = 'b111011000;assign rom[5120] = 'b111011000;assign rom[5121] = 'b101111000;assign rom[5122] = 'b000110011;assign rom[5123] = 'b110000010;assign rom[5124] = 'b001101010;assign rom[5125] = 'b001011000;assign rom[5126] = 'b101001000;assign rom[5127] = 'b000101011;assign rom[5128] = 'b110000010;assign rom[5129] = 'b111000000;assign rom[5130] = 'b101001100;assign rom[5131] = 'b001001010;assign rom[5132] = 'b111111000;assign rom[5133] = 'b111101000;assign rom[5134] = 'b101001111;assign rom[5135] = 'b000111010;assign rom[5136] = 'b101110110;assign rom[5137] = 'b101100010;assign rom[5138] = 'b101001100;assign rom[5139] = 'b001001010;assign rom[5140] = 'b111011010;assign rom[5141] = 'b111011010;assign rom[5142] = 'b111011010;assign rom[5143] = 'b111011010;assign rom[5144] = 'b111011000;assign rom[5145] = 'b111011000;assign rom[5146] = 'b111011000;assign rom[5147] = 'b111011000;assign rom[5148] = 'b101111000;assign rom[5149] = 'b000110011;assign rom[5150] = 'b110000010;assign rom[5151] = 'b001101010;assign rom[5152] = 'b001011000;assign rom[5153] = 'b101001000;assign rom[5154] = 'b000101011;assign rom[5155] = 'b110000010;assign rom[5156] = 'b111000000;assign rom[5157] = 'b101001100;assign rom[5158] = 'b001001010;assign rom[5159] = 'b111111000;assign rom[5160] = 'b111101000;assign rom[5161] = 'b101001111;assign rom[5162] = 'b000111010;assign rom[5163] = 'b101110110;assign rom[5164] = 'b101100010;assign rom[5165] = 'b101001100;assign rom[5166] = 'b001001010;assign rom[5167] = 'b111011010;assign rom[5168] = 'b111011010;assign rom[5169] = 'b111011010;assign rom[5170] = 'b111011010;assign rom[5171] = 'b111011000;assign rom[5172] = 'b111011000;assign rom[5173] = 'b111011000;assign rom[5174] = 'b111011000;assign rom[5175] = 'b101111000;assign rom[5176] = 'b000110011;assign rom[5177] = 'b110000010;assign rom[5178] = 'b001101010;assign rom[5179] = 'b001011000;assign rom[5180] = 'b101001000;assign rom[5181] = 'b000101011;assign rom[5182] = 'b110000010;assign rom[5183] = 'b111000000;assign rom[5184] = 'b101001100;assign rom[5185] = 'b001001010;assign rom[5186] = 'b111111000;assign rom[5187] = 'b111101000;assign rom[5188] = 'b101001111;assign rom[5189] = 'b000111010;assign rom[5190] = 'b101110110;assign rom[5191] = 'b101100010;assign rom[5192] = 'b101001100;assign rom[5193] = 'b001001010;assign rom[5194] = 'b111011010;assign rom[5195] = 'b111011010;assign rom[5196] = 'b111011010;assign rom[5197] = 'b111011010;assign rom[5198] = 'b111011000;assign rom[5199] = 'b111011000;assign rom[5200] = 'b111011000;assign rom[5201] = 'b111011000;assign rom[5202] = 'b101111000;assign rom[5203] = 'b000110011;assign rom[5204] = 'b110000010;assign rom[5205] = 'b001101010;assign rom[5206] = 'b001011000;assign rom[5207] = 'b101001000;assign rom[5208] = 'b000101011;assign rom[5209] = 'b110000010;assign rom[5210] = 'b111000000;assign rom[5211] = 'b101001100;assign rom[5212] = 'b001001010;assign rom[5213] = 'b111111000;assign rom[5214] = 'b111101000;assign rom[5215] = 'b101001111;assign rom[5216] = 'b000111010;assign rom[5217] = 'b101110110;assign rom[5218] = 'b101100010;assign rom[5219] = 'b101001100;assign rom[5220] = 'b001001010;assign rom[5221] = 'b111011010;assign rom[5222] = 'b111011010;assign rom[5223] = 'b111011010;assign rom[5224] = 'b111011010;assign rom[5225] = 'b111011000;assign rom[5226] = 'b111011000;assign rom[5227] = 'b111011000;assign rom[5228] = 'b111011000;assign rom[5229] = 'b101111000;assign rom[5230] = 'b000110011;assign rom[5231] = 'b110000010;assign rom[5232] = 'b001101010;assign rom[5233] = 'b001011000;assign rom[5234] = 'b101001000;assign rom[5235] = 'b000101011;assign rom[5236] = 'b110000010;assign rom[5237] = 'b111000000;assign rom[5238] = 'b101001100;assign rom[5239] = 'b001001010;assign rom[5240] = 'b111111000;assign rom[5241] = 'b111101000;assign rom[5242] = 'b101001111;assign rom[5243] = 'b000111010;assign rom[5244] = 'b101110110;assign rom[5245] = 'b101100010;assign rom[5246] = 'b101001100;assign rom[5247] = 'b001001010;assign rom[5248] = 'b111011010;assign rom[5249] = 'b111011010;assign rom[5250] = 'b111011010;assign rom[5251] = 'b111011010;assign rom[5252] = 'b111011000;assign rom[5253] = 'b111011000;assign rom[5254] = 'b111011000;assign rom[5255] = 'b111011000;assign rom[5256] = 'b101111000;assign rom[5257] = 'b000110011;assign rom[5258] = 'b110000010;assign rom[5259] = 'b001101010;assign rom[5260] = 'b001011000;assign rom[5261] = 'b101001000;assign rom[5262] = 'b000101011;assign rom[5263] = 'b110000010;assign rom[5264] = 'b111000000;assign rom[5265] = 'b101001100;assign rom[5266] = 'b001001010;assign rom[5267] = 'b111111000;assign rom[5268] = 'b111101000;assign rom[5269] = 'b101001111;assign rom[5270] = 'b000111010;assign rom[5271] = 'b101110110;assign rom[5272] = 'b101100010;assign rom[5273] = 'b101001100;assign rom[5274] = 'b001001010;assign rom[5275] = 'b111011010;assign rom[5276] = 'b111011010;assign rom[5277] = 'b111011010;assign rom[5278] = 'b111011010;assign rom[5279] = 'b111011000;assign rom[5280] = 'b111011000;assign rom[5281] = 'b111011000;assign rom[5282] = 'b111011000;assign rom[5283] = 'b101111000;assign rom[5284] = 'b000110011;assign rom[5285] = 'b110000010;assign rom[5286] = 'b001101010;assign rom[5287] = 'b001011000;assign rom[5288] = 'b101001000;assign rom[5289] = 'b000101011;assign rom[5290] = 'b110000010;assign rom[5291] = 'b111000000;assign rom[5292] = 'b101001100;assign rom[5293] = 'b001001010;assign rom[5294] = 'b111111000;assign rom[5295] = 'b111101000;assign rom[5296] = 'b101001111;assign rom[5297] = 'b000111010;assign rom[5298] = 'b101110110;assign rom[5299] = 'b101100010;assign rom[5300] = 'b101001100;assign rom[5301] = 'b001001010;assign rom[5302] = 'b111011010;assign rom[5303] = 'b111011010;assign rom[5304] = 'b111011010;assign rom[5305] = 'b111011010;assign rom[5306] = 'b111011000;assign rom[5307] = 'b111011000;assign rom[5308] = 'b111011000;assign rom[5309] = 'b111011000;assign rom[5310] = 'b101111000;assign rom[5311] = 'b000110011;assign rom[5312] = 'b110000010;assign rom[5313] = 'b001101010;assign rom[5314] = 'b001011000;assign rom[5315] = 'b101001000;assign rom[5316] = 'b000101011;assign rom[5317] = 'b110000010;assign rom[5318] = 'b111000000;assign rom[5319] = 'b101001100;assign rom[5320] = 'b001001010;assign rom[5321] = 'b001000110;assign rom[5322] = 'b001100100;assign rom[5323] = 'b101100010;assign rom[5324] = 'b101001100;assign rom[5325] = 'b001001010;assign rom[5326] = 'b111011010;assign rom[5327] = 'b111011010;assign rom[5328] = 'b111011010;assign rom[5329] = 'b111011010;assign rom[5330] = 'b111011000;assign rom[5331] = 'b111011000;assign rom[5332] = 'b111011000;assign rom[5333] = 'b111011000;assign rom[5334] = 'b101111000;assign rom[5335] = 'b000110011;assign rom[5336] = 'b110000010;assign rom[5337] = 'b001101010;assign rom[5338] = 'b001011000;assign rom[5339] = 'b101001000;assign rom[5340] = 'b000101011;assign rom[5341] = 'b110000010;assign rom[5342] = 'b111000000;assign rom[5343] = 'b101001100;assign rom[5344] = 'b001001010;assign rom[5345] = 'b111111000;assign rom[5346] = 'b111101000;assign rom[5347] = 'b101001111;assign rom[5348] = 'b000111010;assign rom[5349] = 'b101110110;assign rom[5350] = 'b101100010;assign rom[5351] = 'b101001100;assign rom[5352] = 'b001001010;assign rom[5353] = 'b111011010;assign rom[5354] = 'b111011010;assign rom[5355] = 'b111011010;assign rom[5356] = 'b111011010;assign rom[5357] = 'b111011000;assign rom[5358] = 'b111011000;assign rom[5359] = 'b111011000;assign rom[5360] = 'b111011000;assign rom[5361] = 'b101111000;assign rom[5362] = 'b000110011;assign rom[5363] = 'b110000010;assign rom[5364] = 'b001101010;assign rom[5365] = 'b001011000;assign rom[5366] = 'b101001000;assign rom[5367] = 'b000101011;assign rom[5368] = 'b110000010;assign rom[5369] = 'b111000000;assign rom[5370] = 'b101001100;assign rom[5371] = 'b001001010;assign rom[5372] = 'b111111000;assign rom[5373] = 'b111101000;assign rom[5374] = 'b101001111;assign rom[5375] = 'b000111010;assign rom[5376] = 'b101110110;assign rom[5377] = 'b101100010;assign rom[5378] = 'b101001100;assign rom[5379] = 'b001001010;assign rom[5380] = 'b111011010;assign rom[5381] = 'b111011010;assign rom[5382] = 'b111011010;assign rom[5383] = 'b111011010;assign rom[5384] = 'b111011000;assign rom[5385] = 'b111011000;assign rom[5386] = 'b111011000;assign rom[5387] = 'b111011000;assign rom[5388] = 'b101111000;assign rom[5389] = 'b000110011;assign rom[5390] = 'b110000010;assign rom[5391] = 'b001101010;assign rom[5392] = 'b001011000;assign rom[5393] = 'b101001000;assign rom[5394] = 'b000101011;assign rom[5395] = 'b110000010;assign rom[5396] = 'b111000000;assign rom[5397] = 'b101001100;assign rom[5398] = 'b001001010;assign rom[5399] = 'b111111000;assign rom[5400] = 'b111101000;assign rom[5401] = 'b101001111;assign rom[5402] = 'b000111010;assign rom[5403] = 'b101110110;assign rom[5404] = 'b101100010;assign rom[5405] = 'b101001100;assign rom[5406] = 'b001001010;assign rom[5407] = 'b111011010;assign rom[5408] = 'b111011010;assign rom[5409] = 'b111011010;assign rom[5410] = 'b111011010;assign rom[5411] = 'b111011000;assign rom[5412] = 'b111011000;assign rom[5413] = 'b111011000;assign rom[5414] = 'b111011000;assign rom[5415] = 'b101111000;assign rom[5416] = 'b000110011;assign rom[5417] = 'b110000010;assign rom[5418] = 'b001101010;assign rom[5419] = 'b001011000;assign rom[5420] = 'b101001000;assign rom[5421] = 'b000101011;assign rom[5422] = 'b110000010;assign rom[5423] = 'b111000000;assign rom[5424] = 'b101001100;assign rom[5425] = 'b001001010;assign rom[5426] = 'b111111000;assign rom[5427] = 'b111101000;assign rom[5428] = 'b101001111;assign rom[5429] = 'b000111010;assign rom[5430] = 'b101110110;assign rom[5431] = 'b101100010;assign rom[5432] = 'b101001100;assign rom[5433] = 'b001001010;assign rom[5434] = 'b111011010;assign rom[5435] = 'b111011010;assign rom[5436] = 'b111011010;assign rom[5437] = 'b111011010;assign rom[5438] = 'b111011000;assign rom[5439] = 'b111011000;assign rom[5440] = 'b111011000;assign rom[5441] = 'b111011000;assign rom[5442] = 'b101111000;assign rom[5443] = 'b000110011;assign rom[5444] = 'b110000010;assign rom[5445] = 'b001101010;assign rom[5446] = 'b001011000;assign rom[5447] = 'b101001000;assign rom[5448] = 'b000101011;assign rom[5449] = 'b110000010;assign rom[5450] = 'b111000000;assign rom[5451] = 'b101001100;assign rom[5452] = 'b001001010;assign rom[5453] = 'b111111000;assign rom[5454] = 'b111101000;assign rom[5455] = 'b101001111;assign rom[5456] = 'b000111010;assign rom[5457] = 'b101110110;assign rom[5458] = 'b101100010;assign rom[5459] = 'b101001100;assign rom[5460] = 'b001001010;assign rom[5461] = 'b111011010;assign rom[5462] = 'b111011010;assign rom[5463] = 'b111011010;assign rom[5464] = 'b111011010;assign rom[5465] = 'b111011000;assign rom[5466] = 'b111011000;assign rom[5467] = 'b111011000;assign rom[5468] = 'b111011000;assign rom[5469] = 'b101111000;assign rom[5470] = 'b000110011;assign rom[5471] = 'b110000010;assign rom[5472] = 'b001101010;assign rom[5473] = 'b001011000;assign rom[5474] = 'b101001000;assign rom[5475] = 'b000101011;assign rom[5476] = 'b110000010;assign rom[5477] = 'b111000000;assign rom[5478] = 'b101001100;assign rom[5479] = 'b001001010;assign rom[5480] = 'b111111000;assign rom[5481] = 'b111101000;assign rom[5482] = 'b101001111;assign rom[5483] = 'b000111010;assign rom[5484] = 'b101110110;assign rom[5485] = 'b101100010;assign rom[5486] = 'b101001100;assign rom[5487] = 'b001001010;assign rom[5488] = 'b111011010;assign rom[5489] = 'b111011010;assign rom[5490] = 'b111011010;assign rom[5491] = 'b111011010;assign rom[5492] = 'b111011000;assign rom[5493] = 'b111011000;assign rom[5494] = 'b111011000;assign rom[5495] = 'b111011000;assign rom[5496] = 'b101111000;assign rom[5497] = 'b000110011;assign rom[5498] = 'b110000010;assign rom[5499] = 'b001101010;assign rom[5500] = 'b001011000;assign rom[5501] = 'b101001000;assign rom[5502] = 'b000101011;assign rom[5503] = 'b110000010;assign rom[5504] = 'b111000000;assign rom[5505] = 'b101001100;assign rom[5506] = 'b001001010;assign rom[5507] = 'b111111000;assign rom[5508] = 'b111101000;assign rom[5509] = 'b101001111;assign rom[5510] = 'b000111010;assign rom[5511] = 'b101110110;assign rom[5512] = 'b101100010;assign rom[5513] = 'b101001100;assign rom[5514] = 'b001001010;assign rom[5515] = 'b111011010;assign rom[5516] = 'b111011010;assign rom[5517] = 'b111011010;assign rom[5518] = 'b111011010;assign rom[5519] = 'b111011000;assign rom[5520] = 'b111011000;assign rom[5521] = 'b111011000;assign rom[5522] = 'b111011000;assign rom[5523] = 'b101111000;assign rom[5524] = 'b000110011;assign rom[5525] = 'b110000010;assign rom[5526] = 'b001101010;assign rom[5527] = 'b001011000;assign rom[5528] = 'b101001000;assign rom[5529] = 'b000101011;assign rom[5530] = 'b110000010;assign rom[5531] = 'b111000000;assign rom[5532] = 'b101001100;assign rom[5533] = 'b001001010;assign rom[5534] = 'b111111000;assign rom[5535] = 'b111101000;assign rom[5536] = 'b101001111;assign rom[5537] = 'b000111010;assign rom[5538] = 'b101110110;assign rom[5539] = 'b101100010;assign rom[5540] = 'b101001100;assign rom[5541] = 'b001001010;assign rom[5542] = 'b111011010;assign rom[5543] = 'b111011010;assign rom[5544] = 'b111011010;assign rom[5545] = 'b111011010;assign rom[5546] = 'b111011000;assign rom[5547] = 'b111011000;assign rom[5548] = 'b111011000;assign rom[5549] = 'b111011000;assign rom[5550] = 'b101111000;assign rom[5551] = 'b000110011;assign rom[5552] = 'b110000010;assign rom[5553] = 'b001101010;assign rom[5554] = 'b001011000;assign rom[5555] = 'b101001000;assign rom[5556] = 'b000101011;assign rom[5557] = 'b110000010;assign rom[5558] = 'b111000000;assign rom[5559] = 'b101001100;assign rom[5560] = 'b001001010;assign rom[5561] = 'b001000110;assign rom[5562] = 'b001100100;assign rom[5563] = 'b101100010;assign rom[5564] = 'b101001100;assign rom[5565] = 'b001001010;assign rom[5566] = 'b111011010;assign rom[5567] = 'b111011010;assign rom[5568] = 'b111011010;assign rom[5569] = 'b111011010;assign rom[5570] = 'b111011000;assign rom[5571] = 'b111011000;assign rom[5572] = 'b111011000;assign rom[5573] = 'b111011000;assign rom[5574] = 'b101111000;assign rom[5575] = 'b000110011;assign rom[5576] = 'b110000010;assign rom[5577] = 'b001101010;assign rom[5578] = 'b001011000;assign rom[5579] = 'b101001000;assign rom[5580] = 'b000101011;assign rom[5581] = 'b110000010;assign rom[5582] = 'b111000000;assign rom[5583] = 'b101001100;assign rom[5584] = 'b001001010;assign rom[5585] = 'b111111000;assign rom[5586] = 'b111101000;assign rom[5587] = 'b101001111;assign rom[5588] = 'b000111010;assign rom[5589] = 'b101110110;assign rom[5590] = 'b101100010;assign rom[5591] = 'b101001100;assign rom[5592] = 'b001001010;assign rom[5593] = 'b111011010;assign rom[5594] = 'b111011010;assign rom[5595] = 'b111011010;assign rom[5596] = 'b111011010;assign rom[5597] = 'b111011000;assign rom[5598] = 'b111011000;assign rom[5599] = 'b111011000;assign rom[5600] = 'b111011000;assign rom[5601] = 'b101111000;assign rom[5602] = 'b000110011;assign rom[5603] = 'b110000010;assign rom[5604] = 'b001101010;assign rom[5605] = 'b001011000;assign rom[5606] = 'b101001000;assign rom[5607] = 'b000101011;assign rom[5608] = 'b110000010;assign rom[5609] = 'b111000000;assign rom[5610] = 'b101001100;assign rom[5611] = 'b001001010;assign rom[5612] = 'b111111000;assign rom[5613] = 'b111101000;assign rom[5614] = 'b101001111;assign rom[5615] = 'b000111010;assign rom[5616] = 'b101110110;assign rom[5617] = 'b101100010;assign rom[5618] = 'b101001100;assign rom[5619] = 'b001001010;assign rom[5620] = 'b111011010;assign rom[5621] = 'b111011010;assign rom[5622] = 'b111011010;assign rom[5623] = 'b111011010;assign rom[5624] = 'b111011000;assign rom[5625] = 'b111011000;assign rom[5626] = 'b111011000;assign rom[5627] = 'b111011000;assign rom[5628] = 'b101111000;assign rom[5629] = 'b000110011;assign rom[5630] = 'b110000010;assign rom[5631] = 'b001101010;assign rom[5632] = 'b001011000;assign rom[5633] = 'b101001000;assign rom[5634] = 'b000101011;assign rom[5635] = 'b110000010;assign rom[5636] = 'b111000000;assign rom[5637] = 'b101001100;assign rom[5638] = 'b001001010;assign rom[5639] = 'b111111000;assign rom[5640] = 'b111101000;assign rom[5641] = 'b101001111;assign rom[5642] = 'b000111010;assign rom[5643] = 'b101110110;assign rom[5644] = 'b101100010;assign rom[5645] = 'b101001100;assign rom[5646] = 'b001001010;assign rom[5647] = 'b111011010;assign rom[5648] = 'b111011010;assign rom[5649] = 'b111011010;assign rom[5650] = 'b111011010;assign rom[5651] = 'b111011000;assign rom[5652] = 'b111011000;assign rom[5653] = 'b111011000;assign rom[5654] = 'b111011000;assign rom[5655] = 'b101111000;assign rom[5656] = 'b000110011;assign rom[5657] = 'b110000010;assign rom[5658] = 'b001101010;assign rom[5659] = 'b001011000;assign rom[5660] = 'b101001000;assign rom[5661] = 'b000101011;assign rom[5662] = 'b110000010;assign rom[5663] = 'b111000000;assign rom[5664] = 'b101001100;assign rom[5665] = 'b001001010;assign rom[5666] = 'b111111000;assign rom[5667] = 'b111101000;assign rom[5668] = 'b101001111;assign rom[5669] = 'b000111010;assign rom[5670] = 'b101110110;assign rom[5671] = 'b101100010;assign rom[5672] = 'b101001100;assign rom[5673] = 'b001001010;assign rom[5674] = 'b111011010;assign rom[5675] = 'b111011010;assign rom[5676] = 'b111011010;assign rom[5677] = 'b111011010;assign rom[5678] = 'b111011000;assign rom[5679] = 'b111011000;assign rom[5680] = 'b111011000;assign rom[5681] = 'b111011000;assign rom[5682] = 'b101111000;assign rom[5683] = 'b000110011;assign rom[5684] = 'b110000010;assign rom[5685] = 'b001101010;assign rom[5686] = 'b001011000;assign rom[5687] = 'b101001000;assign rom[5688] = 'b000101011;assign rom[5689] = 'b110000010;assign rom[5690] = 'b111000000;assign rom[5691] = 'b101001100;assign rom[5692] = 'b001001010;assign rom[5693] = 'b111111000;assign rom[5694] = 'b111101000;assign rom[5695] = 'b101001111;assign rom[5696] = 'b000111010;assign rom[5697] = 'b101110110;assign rom[5698] = 'b101100010;assign rom[5699] = 'b101001100;assign rom[5700] = 'b001001010;assign rom[5701] = 'b111011010;assign rom[5702] = 'b111011010;assign rom[5703] = 'b111011010;assign rom[5704] = 'b111011010;assign rom[5705] = 'b111011000;assign rom[5706] = 'b111011000;assign rom[5707] = 'b111011000;assign rom[5708] = 'b111011000;assign rom[5709] = 'b101111000;assign rom[5710] = 'b000110011;assign rom[5711] = 'b110000010;assign rom[5712] = 'b001101010;assign rom[5713] = 'b001011000;assign rom[5714] = 'b101001000;assign rom[5715] = 'b000101011;assign rom[5716] = 'b110000010;assign rom[5717] = 'b111000000;assign rom[5718] = 'b101001100;assign rom[5719] = 'b001001010;assign rom[5720] = 'b111111000;assign rom[5721] = 'b111101000;assign rom[5722] = 'b101001111;assign rom[5723] = 'b000111010;assign rom[5724] = 'b101110110;assign rom[5725] = 'b101100010;assign rom[5726] = 'b101001100;assign rom[5727] = 'b001001010;assign rom[5728] = 'b111011010;assign rom[5729] = 'b111011010;assign rom[5730] = 'b111011010;assign rom[5731] = 'b111011010;assign rom[5732] = 'b111011000;assign rom[5733] = 'b111011000;assign rom[5734] = 'b111011000;assign rom[5735] = 'b111011000;assign rom[5736] = 'b101111000;assign rom[5737] = 'b000110011;assign rom[5738] = 'b110000010;assign rom[5739] = 'b001101010;assign rom[5740] = 'b001011000;assign rom[5741] = 'b101001000;assign rom[5742] = 'b000101011;assign rom[5743] = 'b110000010;assign rom[5744] = 'b111000000;assign rom[5745] = 'b101001100;assign rom[5746] = 'b001001010;assign rom[5747] = 'b111111000;assign rom[5748] = 'b111101000;assign rom[5749] = 'b101001111;assign rom[5750] = 'b000111010;assign rom[5751] = 'b101110110;assign rom[5752] = 'b101100010;assign rom[5753] = 'b101001100;assign rom[5754] = 'b001001010;assign rom[5755] = 'b111011010;assign rom[5756] = 'b111011010;assign rom[5757] = 'b111011010;assign rom[5758] = 'b111011010;assign rom[5759] = 'b111011000;assign rom[5760] = 'b111011000;assign rom[5761] = 'b111011000;assign rom[5762] = 'b111011000;assign rom[5763] = 'b101111000;assign rom[5764] = 'b000110011;assign rom[5765] = 'b110000010;assign rom[5766] = 'b001101010;assign rom[5767] = 'b001011000;assign rom[5768] = 'b101001000;assign rom[5769] = 'b000101011;assign rom[5770] = 'b110000010;assign rom[5771] = 'b111000000;assign rom[5772] = 'b101001100;assign rom[5773] = 'b001001010;assign rom[5774] = 'b111111000;assign rom[5775] = 'b111101000;assign rom[5776] = 'b101001111;assign rom[5777] = 'b000111010;assign rom[5778] = 'b101110110;assign rom[5779] = 'b101100010;assign rom[5780] = 'b101001100;assign rom[5781] = 'b001001010;assign rom[5782] = 'b111011010;assign rom[5783] = 'b111011010;assign rom[5784] = 'b111011010;assign rom[5785] = 'b111011010;assign rom[5786] = 'b111011000;assign rom[5787] = 'b111011000;assign rom[5788] = 'b111011000;assign rom[5789] = 'b111011000;assign rom[5790] = 'b101111000;assign rom[5791] = 'b000110011;assign rom[5792] = 'b110000010;assign rom[5793] = 'b001101010;assign rom[5794] = 'b001011000;assign rom[5795] = 'b101001000;assign rom[5796] = 'b000101011;assign rom[5797] = 'b110000010;assign rom[5798] = 'b111000000;assign rom[5799] = 'b101001100;assign rom[5800] = 'b001001010;assign rom[5801] = 'b001000110;assign rom[5802] = 'b001100100;assign rom[5803] = 'b101100010;assign rom[5804] = 'b101001100;assign rom[5805] = 'b001001010;assign rom[5806] = 'b111011010;assign rom[5807] = 'b111011010;assign rom[5808] = 'b111011010;assign rom[5809] = 'b111011010;assign rom[5810] = 'b111011000;assign rom[5811] = 'b111011000;assign rom[5812] = 'b111011000;assign rom[5813] = 'b111011000;assign rom[5814] = 'b101111000;assign rom[5815] = 'b000110011;assign rom[5816] = 'b110000010;assign rom[5817] = 'b001101010;assign rom[5818] = 'b001011000;assign rom[5819] = 'b101001000;assign rom[5820] = 'b000101011;assign rom[5821] = 'b110000010;assign rom[5822] = 'b111000000;assign rom[5823] = 'b101001100;assign rom[5824] = 'b001001010;assign rom[5825] = 'b111111000;assign rom[5826] = 'b111101000;assign rom[5827] = 'b101001111;assign rom[5828] = 'b000111010;assign rom[5829] = 'b101110110;assign rom[5830] = 'b101100010;assign rom[5831] = 'b101001100;assign rom[5832] = 'b001001010;assign rom[5833] = 'b111011010;assign rom[5834] = 'b111011010;assign rom[5835] = 'b111011010;assign rom[5836] = 'b111011010;assign rom[5837] = 'b111011000;assign rom[5838] = 'b111011000;assign rom[5839] = 'b111011000;assign rom[5840] = 'b111011000;assign rom[5841] = 'b101111000;assign rom[5842] = 'b000110011;assign rom[5843] = 'b110000010;assign rom[5844] = 'b001101010;assign rom[5845] = 'b001011000;assign rom[5846] = 'b101001000;assign rom[5847] = 'b000101011;assign rom[5848] = 'b110000010;assign rom[5849] = 'b111000000;assign rom[5850] = 'b101001100;assign rom[5851] = 'b001001010;assign rom[5852] = 'b111111000;assign rom[5853] = 'b111101000;assign rom[5854] = 'b101001111;assign rom[5855] = 'b000111010;assign rom[5856] = 'b101110110;assign rom[5857] = 'b101100010;assign rom[5858] = 'b101001100;assign rom[5859] = 'b001001010;assign rom[5860] = 'b111011010;assign rom[5861] = 'b111011010;assign rom[5862] = 'b111011010;assign rom[5863] = 'b111011010;assign rom[5864] = 'b111011000;assign rom[5865] = 'b111011000;assign rom[5866] = 'b111011000;assign rom[5867] = 'b111011000;assign rom[5868] = 'b101111000;assign rom[5869] = 'b000110011;assign rom[5870] = 'b110000010;assign rom[5871] = 'b001101010;assign rom[5872] = 'b001011000;assign rom[5873] = 'b101001000;assign rom[5874] = 'b000101011;assign rom[5875] = 'b110000010;assign rom[5876] = 'b111000000;assign rom[5877] = 'b101001100;assign rom[5878] = 'b001001010;assign rom[5879] = 'b111111000;assign rom[5880] = 'b111101000;assign rom[5881] = 'b101001111;assign rom[5882] = 'b000111010;assign rom[5883] = 'b101110110;assign rom[5884] = 'b101100010;assign rom[5885] = 'b101001100;assign rom[5886] = 'b001001010;assign rom[5887] = 'b111011010;assign rom[5888] = 'b111011010;assign rom[5889] = 'b111011010;assign rom[5890] = 'b111011010;assign rom[5891] = 'b111011000;assign rom[5892] = 'b111011000;assign rom[5893] = 'b111011000;assign rom[5894] = 'b111011000;assign rom[5895] = 'b101111000;assign rom[5896] = 'b000110011;assign rom[5897] = 'b110000010;assign rom[5898] = 'b001101010;assign rom[5899] = 'b001011000;assign rom[5900] = 'b101001000;assign rom[5901] = 'b000101011;assign rom[5902] = 'b110000010;assign rom[5903] = 'b111000000;assign rom[5904] = 'b101001100;assign rom[5905] = 'b001001010;assign rom[5906] = 'b111111000;assign rom[5907] = 'b111101000;assign rom[5908] = 'b101001111;assign rom[5909] = 'b000111010;assign rom[5910] = 'b101110110;assign rom[5911] = 'b101100010;assign rom[5912] = 'b101001100;assign rom[5913] = 'b001001010;assign rom[5914] = 'b111011010;assign rom[5915] = 'b111011010;assign rom[5916] = 'b111011010;assign rom[5917] = 'b111011010;assign rom[5918] = 'b111011000;assign rom[5919] = 'b111011000;assign rom[5920] = 'b111011000;assign rom[5921] = 'b111011000;assign rom[5922] = 'b101111000;assign rom[5923] = 'b000110011;assign rom[5924] = 'b110000010;assign rom[5925] = 'b001101010;assign rom[5926] = 'b001011000;assign rom[5927] = 'b101001000;assign rom[5928] = 'b000101011;assign rom[5929] = 'b110000010;assign rom[5930] = 'b111000000;assign rom[5931] = 'b101001100;assign rom[5932] = 'b001001010;assign rom[5933] = 'b111111000;assign rom[5934] = 'b111101000;assign rom[5935] = 'b101001111;assign rom[5936] = 'b000111010;assign rom[5937] = 'b101110110;assign rom[5938] = 'b101100010;assign rom[5939] = 'b101001100;assign rom[5940] = 'b001001010;assign rom[5941] = 'b111011010;assign rom[5942] = 'b111011010;assign rom[5943] = 'b111011010;assign rom[5944] = 'b111011010;assign rom[5945] = 'b111011000;assign rom[5946] = 'b111011000;assign rom[5947] = 'b111011000;assign rom[5948] = 'b111011000;assign rom[5949] = 'b101111000;assign rom[5950] = 'b000110011;assign rom[5951] = 'b110000010;assign rom[5952] = 'b001101010;assign rom[5953] = 'b001011000;assign rom[5954] = 'b101001000;assign rom[5955] = 'b000101011;assign rom[5956] = 'b110000010;assign rom[5957] = 'b111000000;assign rom[5958] = 'b101001100;assign rom[5959] = 'b001001010;assign rom[5960] = 'b111111000;assign rom[5961] = 'b111101000;assign rom[5962] = 'b101001111;assign rom[5963] = 'b000111010;assign rom[5964] = 'b101110110;assign rom[5965] = 'b101100010;assign rom[5966] = 'b101001100;assign rom[5967] = 'b001001010;assign rom[5968] = 'b111011010;assign rom[5969] = 'b111011010;assign rom[5970] = 'b111011010;assign rom[5971] = 'b111011010;assign rom[5972] = 'b111011000;assign rom[5973] = 'b111011000;assign rom[5974] = 'b111011000;assign rom[5975] = 'b111011000;assign rom[5976] = 'b101111000;assign rom[5977] = 'b000110011;assign rom[5978] = 'b110000010;assign rom[5979] = 'b001101010;assign rom[5980] = 'b001011000;assign rom[5981] = 'b101001000;assign rom[5982] = 'b000101011;assign rom[5983] = 'b110000010;assign rom[5984] = 'b111000000;assign rom[5985] = 'b101001100;assign rom[5986] = 'b001001010;assign rom[5987] = 'b111111000;assign rom[5988] = 'b111101000;assign rom[5989] = 'b101001111;assign rom[5990] = 'b000111010;assign rom[5991] = 'b101110110;assign rom[5992] = 'b101100010;assign rom[5993] = 'b101001100;assign rom[5994] = 'b001001010;assign rom[5995] = 'b111011010;assign rom[5996] = 'b111011010;assign rom[5997] = 'b111011010;assign rom[5998] = 'b111011010;assign rom[5999] = 'b111011000;assign rom[6000] = 'b111011000;assign rom[6001] = 'b111011000;assign rom[6002] = 'b111011000;assign rom[6003] = 'b101111000;assign rom[6004] = 'b000110011;assign rom[6005] = 'b110000010;assign rom[6006] = 'b001101010;assign rom[6007] = 'b001011000;assign rom[6008] = 'b101001000;assign rom[6009] = 'b000101011;assign rom[6010] = 'b110000010;assign rom[6011] = 'b111000000;assign rom[6012] = 'b101001100;assign rom[6013] = 'b001001010;assign rom[6014] = 'b111111000;assign rom[6015] = 'b111101000;assign rom[6016] = 'b101001111;assign rom[6017] = 'b000111010;assign rom[6018] = 'b101110110;assign rom[6019] = 'b101100010;assign rom[6020] = 'b101001100;assign rom[6021] = 'b001001010;assign rom[6022] = 'b111011010;assign rom[6023] = 'b111011010;assign rom[6024] = 'b111011010;assign rom[6025] = 'b111011010;assign rom[6026] = 'b111011000;assign rom[6027] = 'b111011000;assign rom[6028] = 'b111011000;assign rom[6029] = 'b111011000;assign rom[6030] = 'b101111000;assign rom[6031] = 'b000110011;assign rom[6032] = 'b110000010;assign rom[6033] = 'b001101010;assign rom[6034] = 'b001011000;assign rom[6035] = 'b101001000;assign rom[6036] = 'b000101011;assign rom[6037] = 'b110000010;assign rom[6038] = 'b111000000;assign rom[6039] = 'b101001100;assign rom[6040] = 'b001001010;assign rom[6041] = 'b001000110;assign rom[6042] = 'b001100100;assign rom[6043] = 'b101100010;assign rom[6044] = 'b101001100;assign rom[6045] = 'b001001010;assign rom[6046] = 'b111011010;assign rom[6047] = 'b111011010;assign rom[6048] = 'b111011010;assign rom[6049] = 'b111011010;assign rom[6050] = 'b111011000;assign rom[6051] = 'b111011000;assign rom[6052] = 'b111011000;assign rom[6053] = 'b111011000;assign rom[6054] = 'b101111000;assign rom[6055] = 'b000110011;assign rom[6056] = 'b110000010;assign rom[6057] = 'b001101010;assign rom[6058] = 'b001011000;assign rom[6059] = 'b101001000;assign rom[6060] = 'b000101011;assign rom[6061] = 'b110000010;assign rom[6062] = 'b111000000;assign rom[6063] = 'b101001100;assign rom[6064] = 'b001001010;assign rom[6065] = 'b111111000;assign rom[6066] = 'b111101000;assign rom[6067] = 'b101001111;assign rom[6068] = 'b000111010;assign rom[6069] = 'b101110110;assign rom[6070] = 'b101100010;assign rom[6071] = 'b101001100;assign rom[6072] = 'b001001010;assign rom[6073] = 'b111011010;assign rom[6074] = 'b111011010;assign rom[6075] = 'b111011010;assign rom[6076] = 'b111011010;assign rom[6077] = 'b111011000;assign rom[6078] = 'b111011000;assign rom[6079] = 'b111011000;assign rom[6080] = 'b111011000;assign rom[6081] = 'b101111000;assign rom[6082] = 'b000110011;assign rom[6083] = 'b110000010;assign rom[6084] = 'b001101010;assign rom[6085] = 'b001011000;assign rom[6086] = 'b101001000;assign rom[6087] = 'b000101011;assign rom[6088] = 'b110000010;assign rom[6089] = 'b111000000;assign rom[6090] = 'b101001100;assign rom[6091] = 'b001001010;assign rom[6092] = 'b111111000;assign rom[6093] = 'b111101000;assign rom[6094] = 'b101001111;assign rom[6095] = 'b000111010;assign rom[6096] = 'b101110110;assign rom[6097] = 'b101100010;assign rom[6098] = 'b101001100;assign rom[6099] = 'b001001010;assign rom[6100] = 'b111011010;assign rom[6101] = 'b111011010;assign rom[6102] = 'b111011010;assign rom[6103] = 'b111011010;assign rom[6104] = 'b111011000;assign rom[6105] = 'b111011000;assign rom[6106] = 'b111011000;assign rom[6107] = 'b111011000;assign rom[6108] = 'b101111000;assign rom[6109] = 'b000110011;assign rom[6110] = 'b110000010;assign rom[6111] = 'b001101010;assign rom[6112] = 'b001011000;assign rom[6113] = 'b101001000;assign rom[6114] = 'b000101011;assign rom[6115] = 'b110000010;assign rom[6116] = 'b111000000;assign rom[6117] = 'b101001100;assign rom[6118] = 'b001001010;assign rom[6119] = 'b111111000;assign rom[6120] = 'b111101000;assign rom[6121] = 'b101001111;assign rom[6122] = 'b000111010;assign rom[6123] = 'b101110110;assign rom[6124] = 'b101100010;assign rom[6125] = 'b101001100;assign rom[6126] = 'b001001010;assign rom[6127] = 'b111011010;assign rom[6128] = 'b111011010;assign rom[6129] = 'b111011010;assign rom[6130] = 'b111011010;assign rom[6131] = 'b111011000;assign rom[6132] = 'b111011000;assign rom[6133] = 'b111011000;assign rom[6134] = 'b111011000;assign rom[6135] = 'b101111000;assign rom[6136] = 'b000110011;assign rom[6137] = 'b110000010;assign rom[6138] = 'b001101010;assign rom[6139] = 'b001011000;assign rom[6140] = 'b101001000;assign rom[6141] = 'b000101011;assign rom[6142] = 'b110000010;assign rom[6143] = 'b111000000;assign rom[6144] = 'b101001100;assign rom[6145] = 'b001001010;assign rom[6146] = 'b111111000;assign rom[6147] = 'b111101000;assign rom[6148] = 'b101001111;assign rom[6149] = 'b000111010;assign rom[6150] = 'b101110110;assign rom[6151] = 'b101100010;assign rom[6152] = 'b101001100;assign rom[6153] = 'b001001010;assign rom[6154] = 'b111011010;assign rom[6155] = 'b111011010;assign rom[6156] = 'b111011010;assign rom[6157] = 'b111011010;assign rom[6158] = 'b111011000;assign rom[6159] = 'b111011000;assign rom[6160] = 'b111011000;assign rom[6161] = 'b111011000;assign rom[6162] = 'b101111000;assign rom[6163] = 'b000110011;assign rom[6164] = 'b110000010;assign rom[6165] = 'b001101010;assign rom[6166] = 'b001011000;assign rom[6167] = 'b101001000;assign rom[6168] = 'b000101011;assign rom[6169] = 'b110000010;assign rom[6170] = 'b111000000;assign rom[6171] = 'b101001100;assign rom[6172] = 'b001001010;assign rom[6173] = 'b111111000;assign rom[6174] = 'b111101000;assign rom[6175] = 'b101001111;assign rom[6176] = 'b000111010;assign rom[6177] = 'b101110110;assign rom[6178] = 'b101100010;assign rom[6179] = 'b101001100;assign rom[6180] = 'b001001010;assign rom[6181] = 'b111011010;assign rom[6182] = 'b111011010;assign rom[6183] = 'b111011010;assign rom[6184] = 'b111011010;assign rom[6185] = 'b111011000;assign rom[6186] = 'b111011000;assign rom[6187] = 'b111011000;assign rom[6188] = 'b111011000;assign rom[6189] = 'b101111000;assign rom[6190] = 'b000110011;assign rom[6191] = 'b110000010;assign rom[6192] = 'b001101010;assign rom[6193] = 'b001011000;assign rom[6194] = 'b101001000;assign rom[6195] = 'b000101011;assign rom[6196] = 'b110000010;assign rom[6197] = 'b111000000;assign rom[6198] = 'b101001100;assign rom[6199] = 'b001001010;assign rom[6200] = 'b111111000;assign rom[6201] = 'b111101000;assign rom[6202] = 'b101001111;assign rom[6203] = 'b000111010;assign rom[6204] = 'b101110110;assign rom[6205] = 'b101100010;assign rom[6206] = 'b101001100;assign rom[6207] = 'b001001010;assign rom[6208] = 'b111011010;assign rom[6209] = 'b111011010;assign rom[6210] = 'b111011010;assign rom[6211] = 'b111011010;assign rom[6212] = 'b111011000;assign rom[6213] = 'b111011000;assign rom[6214] = 'b111011000;assign rom[6215] = 'b111011000;assign rom[6216] = 'b101111000;assign rom[6217] = 'b000110011;assign rom[6218] = 'b110000010;assign rom[6219] = 'b001101010;assign rom[6220] = 'b001011000;assign rom[6221] = 'b101001000;assign rom[6222] = 'b000101011;assign rom[6223] = 'b110000010;assign rom[6224] = 'b111000000;assign rom[6225] = 'b101001100;assign rom[6226] = 'b001001010;assign rom[6227] = 'b111111000;assign rom[6228] = 'b111101000;assign rom[6229] = 'b101001111;assign rom[6230] = 'b000111010;assign rom[6231] = 'b101110110;assign rom[6232] = 'b101100010;assign rom[6233] = 'b101001100;assign rom[6234] = 'b001001010;assign rom[6235] = 'b111011010;assign rom[6236] = 'b111011010;assign rom[6237] = 'b111011010;assign rom[6238] = 'b111011010;assign rom[6239] = 'b111011000;assign rom[6240] = 'b111011000;assign rom[6241] = 'b111011000;assign rom[6242] = 'b111011000;assign rom[6243] = 'b101111000;assign rom[6244] = 'b000110011;assign rom[6245] = 'b110000010;assign rom[6246] = 'b001101010;assign rom[6247] = 'b001011000;assign rom[6248] = 'b101001000;assign rom[6249] = 'b000101011;assign rom[6250] = 'b110000010;assign rom[6251] = 'b111000000;assign rom[6252] = 'b101001100;assign rom[6253] = 'b001001010;assign rom[6254] = 'b111111000;assign rom[6255] = 'b111101000;assign rom[6256] = 'b101001111;assign rom[6257] = 'b000111010;assign rom[6258] = 'b101110110;assign rom[6259] = 'b101100010;assign rom[6260] = 'b101001100;assign rom[6261] = 'b001001010;assign rom[6262] = 'b111011010;assign rom[6263] = 'b111011010;assign rom[6264] = 'b111011010;assign rom[6265] = 'b111011010;assign rom[6266] = 'b111011000;assign rom[6267] = 'b111011000;assign rom[6268] = 'b111011000;assign rom[6269] = 'b111011000;assign rom[6270] = 'b101111000;assign rom[6271] = 'b000110011;assign rom[6272] = 'b110000010;assign rom[6273] = 'b001101010;assign rom[6274] = 'b001011000;assign rom[6275] = 'b101001000;assign rom[6276] = 'b000101011;assign rom[6277] = 'b110000010;assign rom[6278] = 'b111000000;assign rom[6279] = 'b101001100;assign rom[6280] = 'b001001010;assign rom[6281] = 'b001000110;assign rom[6282] = 'b001100100;assign rom[6283] = 'b101100010;assign rom[6284] = 'b101001100;assign rom[6285] = 'b001001010;assign rom[6286] = 'b111011010;assign rom[6287] = 'b111011010;assign rom[6288] = 'b111011010;assign rom[6289] = 'b111011010;assign rom[6290] = 'b111011000;assign rom[6291] = 'b111011000;assign rom[6292] = 'b111011000;assign rom[6293] = 'b111011000;assign rom[6294] = 'b101111000;assign rom[6295] = 'b000110011;assign rom[6296] = 'b110000010;assign rom[6297] = 'b001101010;assign rom[6298] = 'b001011000;assign rom[6299] = 'b101001000;assign rom[6300] = 'b000101011;assign rom[6301] = 'b110000010;assign rom[6302] = 'b111000000;assign rom[6303] = 'b101001100;assign rom[6304] = 'b001001010;assign rom[6305] = 'b111111000;assign rom[6306] = 'b111101000;assign rom[6307] = 'b101001111;assign rom[6308] = 'b000111010;assign rom[6309] = 'b101110110;assign rom[6310] = 'b101100010;assign rom[6311] = 'b101001100;assign rom[6312] = 'b001001010;assign rom[6313] = 'b111011010;assign rom[6314] = 'b111011010;assign rom[6315] = 'b111011010;assign rom[6316] = 'b111011010;assign rom[6317] = 'b111011000;assign rom[6318] = 'b111011000;assign rom[6319] = 'b111011000;assign rom[6320] = 'b111011000;assign rom[6321] = 'b101111000;assign rom[6322] = 'b000110011;assign rom[6323] = 'b110000010;assign rom[6324] = 'b001101010;assign rom[6325] = 'b001011000;assign rom[6326] = 'b101001000;assign rom[6327] = 'b000101011;assign rom[6328] = 'b110000010;assign rom[6329] = 'b111000000;assign rom[6330] = 'b101001100;assign rom[6331] = 'b001001010;assign rom[6332] = 'b111111000;assign rom[6333] = 'b111101000;assign rom[6334] = 'b101001111;assign rom[6335] = 'b000111010;assign rom[6336] = 'b101110110;assign rom[6337] = 'b101100010;assign rom[6338] = 'b101001100;assign rom[6339] = 'b001001010;assign rom[6340] = 'b111011010;assign rom[6341] = 'b111011010;assign rom[6342] = 'b111011010;assign rom[6343] = 'b111011010;assign rom[6344] = 'b111011000;assign rom[6345] = 'b111011000;assign rom[6346] = 'b111011000;assign rom[6347] = 'b111011000;assign rom[6348] = 'b101111000;assign rom[6349] = 'b000110011;assign rom[6350] = 'b110000010;assign rom[6351] = 'b001101010;assign rom[6352] = 'b001011000;assign rom[6353] = 'b101001000;assign rom[6354] = 'b000101011;assign rom[6355] = 'b110000010;assign rom[6356] = 'b111000000;assign rom[6357] = 'b101001100;assign rom[6358] = 'b001001010;assign rom[6359] = 'b111111000;assign rom[6360] = 'b111101000;assign rom[6361] = 'b101001111;assign rom[6362] = 'b000111010;assign rom[6363] = 'b101110110;assign rom[6364] = 'b101100010;assign rom[6365] = 'b101001100;assign rom[6366] = 'b001001010;assign rom[6367] = 'b111011010;assign rom[6368] = 'b111011010;assign rom[6369] = 'b111011010;assign rom[6370] = 'b111011010;assign rom[6371] = 'b111011000;assign rom[6372] = 'b111011000;assign rom[6373] = 'b111011000;assign rom[6374] = 'b111011000;assign rom[6375] = 'b101111000;assign rom[6376] = 'b000110011;assign rom[6377] = 'b110000010;assign rom[6378] = 'b001101010;assign rom[6379] = 'b001011000;assign rom[6380] = 'b101001000;assign rom[6381] = 'b000101011;assign rom[6382] = 'b110000010;assign rom[6383] = 'b111000000;assign rom[6384] = 'b101001100;assign rom[6385] = 'b001001010;assign rom[6386] = 'b111111000;assign rom[6387] = 'b111101000;assign rom[6388] = 'b101001111;assign rom[6389] = 'b000111010;assign rom[6390] = 'b101110110;assign rom[6391] = 'b101100010;assign rom[6392] = 'b101001100;assign rom[6393] = 'b001001010;assign rom[6394] = 'b111011010;assign rom[6395] = 'b111011010;assign rom[6396] = 'b111011010;assign rom[6397] = 'b111011010;assign rom[6398] = 'b111011000;assign rom[6399] = 'b111011000;assign rom[6400] = 'b111011000;assign rom[6401] = 'b111011000;assign rom[6402] = 'b101111000;assign rom[6403] = 'b000110011;assign rom[6404] = 'b110000010;assign rom[6405] = 'b001101010;assign rom[6406] = 'b001011000;assign rom[6407] = 'b101001000;assign rom[6408] = 'b000101011;assign rom[6409] = 'b110000010;assign rom[6410] = 'b111000000;assign rom[6411] = 'b101001100;assign rom[6412] = 'b001001010;assign rom[6413] = 'b111111000;assign rom[6414] = 'b111101000;assign rom[6415] = 'b101001111;assign rom[6416] = 'b000111010;assign rom[6417] = 'b101110110;assign rom[6418] = 'b101100010;assign rom[6419] = 'b101001100;assign rom[6420] = 'b001001010;assign rom[6421] = 'b111011010;assign rom[6422] = 'b111011010;assign rom[6423] = 'b111011010;assign rom[6424] = 'b111011010;assign rom[6425] = 'b111011000;assign rom[6426] = 'b111011000;assign rom[6427] = 'b111011000;assign rom[6428] = 'b111011000;assign rom[6429] = 'b101111000;assign rom[6430] = 'b000110011;assign rom[6431] = 'b110000010;assign rom[6432] = 'b001101010;assign rom[6433] = 'b001011000;assign rom[6434] = 'b101001000;assign rom[6435] = 'b000101011;assign rom[6436] = 'b110000010;assign rom[6437] = 'b111000000;assign rom[6438] = 'b101001100;assign rom[6439] = 'b001001010;assign rom[6440] = 'b111111000;assign rom[6441] = 'b111101000;assign rom[6442] = 'b101001111;assign rom[6443] = 'b000111010;assign rom[6444] = 'b101110110;assign rom[6445] = 'b101100010;assign rom[6446] = 'b101001100;assign rom[6447] = 'b001001010;assign rom[6448] = 'b111011010;assign rom[6449] = 'b111011010;assign rom[6450] = 'b111011010;assign rom[6451] = 'b111011010;assign rom[6452] = 'b111011000;assign rom[6453] = 'b111011000;assign rom[6454] = 'b111011000;assign rom[6455] = 'b111011000;assign rom[6456] = 'b101111000;assign rom[6457] = 'b000110011;assign rom[6458] = 'b110000010;assign rom[6459] = 'b001101010;assign rom[6460] = 'b001011000;assign rom[6461] = 'b101001000;assign rom[6462] = 'b000101011;assign rom[6463] = 'b110000010;assign rom[6464] = 'b111000000;assign rom[6465] = 'b101001100;assign rom[6466] = 'b001001010;assign rom[6467] = 'b111111000;assign rom[6468] = 'b111101000;assign rom[6469] = 'b101001111;assign rom[6470] = 'b000111010;assign rom[6471] = 'b101110110;assign rom[6472] = 'b101100010;assign rom[6473] = 'b101001100;assign rom[6474] = 'b001001010;assign rom[6475] = 'b111011010;assign rom[6476] = 'b111011010;assign rom[6477] = 'b111011010;assign rom[6478] = 'b111011010;assign rom[6479] = 'b111011000;assign rom[6480] = 'b111011000;assign rom[6481] = 'b111011000;assign rom[6482] = 'b111011000;assign rom[6483] = 'b101111000;assign rom[6484] = 'b000110011;assign rom[6485] = 'b110000010;assign rom[6486] = 'b001101010;assign rom[6487] = 'b001011000;assign rom[6488] = 'b101001000;assign rom[6489] = 'b000101011;assign rom[6490] = 'b110000010;assign rom[6491] = 'b111000000;assign rom[6492] = 'b101001100;assign rom[6493] = 'b001001010;assign rom[6494] = 'b111111000;assign rom[6495] = 'b111101000;assign rom[6496] = 'b101001111;assign rom[6497] = 'b000111010;assign rom[6498] = 'b101110110;assign rom[6499] = 'b101100010;assign rom[6500] = 'b101001100;assign rom[6501] = 'b001001010;assign rom[6502] = 'b111011010;assign rom[6503] = 'b111011010;assign rom[6504] = 'b111011010;assign rom[6505] = 'b111011010;assign rom[6506] = 'b111011000;assign rom[6507] = 'b111011000;assign rom[6508] = 'b111011000;assign rom[6509] = 'b111011000;assign rom[6510] = 'b101111000;assign rom[6511] = 'b000110011;assign rom[6512] = 'b110000010;assign rom[6513] = 'b001101010;assign rom[6514] = 'b001011000;assign rom[6515] = 'b101001000;assign rom[6516] = 'b000101011;assign rom[6517] = 'b110000010;assign rom[6518] = 'b111000000;assign rom[6519] = 'b101001100;assign rom[6520] = 'b001001010;assign rom[6521] = 'b001000110;assign rom[6522] = 'b001100100;assign rom[6523] = 'b101100010;assign rom[6524] = 'b101001100;assign rom[6525] = 'b001001010;assign rom[6526] = 'b111011010;assign rom[6527] = 'b111011010;assign rom[6528] = 'b111011010;assign rom[6529] = 'b111011010;assign rom[6530] = 'b111011000;assign rom[6531] = 'b111011000;assign rom[6532] = 'b111011000;assign rom[6533] = 'b111011000;assign rom[6534] = 'b101111000;assign rom[6535] = 'b000110011;assign rom[6536] = 'b110000010;assign rom[6537] = 'b001101010;assign rom[6538] = 'b001011000;assign rom[6539] = 'b101001000;assign rom[6540] = 'b000101011;assign rom[6541] = 'b110000010;assign rom[6542] = 'b111000000;assign rom[6543] = 'b101001100;assign rom[6544] = 'b001001010;assign rom[6545] = 'b111111000;assign rom[6546] = 'b111101000;assign rom[6547] = 'b101001111;assign rom[6548] = 'b000111010;assign rom[6549] = 'b101110110;assign rom[6550] = 'b101100010;assign rom[6551] = 'b101001100;assign rom[6552] = 'b001001010;assign rom[6553] = 'b111011010;assign rom[6554] = 'b111011010;assign rom[6555] = 'b111011010;assign rom[6556] = 'b111011010;assign rom[6557] = 'b111011000;assign rom[6558] = 'b111011000;assign rom[6559] = 'b111011000;assign rom[6560] = 'b111011000;assign rom[6561] = 'b101111000;assign rom[6562] = 'b000110011;assign rom[6563] = 'b110000010;assign rom[6564] = 'b001101010;assign rom[6565] = 'b001011000;assign rom[6566] = 'b101001000;assign rom[6567] = 'b000101011;assign rom[6568] = 'b110000010;assign rom[6569] = 'b111000000;assign rom[6570] = 'b101001100;assign rom[6571] = 'b001001010;assign rom[6572] = 'b111111000;assign rom[6573] = 'b111101000;assign rom[6574] = 'b101001111;assign rom[6575] = 'b000111010;assign rom[6576] = 'b101110110;assign rom[6577] = 'b101100010;assign rom[6578] = 'b101001100;assign rom[6579] = 'b001001010;assign rom[6580] = 'b111011010;assign rom[6581] = 'b111011010;assign rom[6582] = 'b111011010;assign rom[6583] = 'b111011010;assign rom[6584] = 'b111011000;assign rom[6585] = 'b111011000;assign rom[6586] = 'b111011000;assign rom[6587] = 'b111011000;assign rom[6588] = 'b101111000;assign rom[6589] = 'b000110011;assign rom[6590] = 'b110000010;assign rom[6591] = 'b001101010;assign rom[6592] = 'b001011000;assign rom[6593] = 'b101001000;assign rom[6594] = 'b000101011;assign rom[6595] = 'b110000010;assign rom[6596] = 'b111000000;assign rom[6597] = 'b101001100;assign rom[6598] = 'b001001010;assign rom[6599] = 'b111111000;assign rom[6600] = 'b111101000;assign rom[6601] = 'b101001111;assign rom[6602] = 'b000111010;assign rom[6603] = 'b101110110;assign rom[6604] = 'b101100010;assign rom[6605] = 'b101001100;assign rom[6606] = 'b001001010;assign rom[6607] = 'b111011010;assign rom[6608] = 'b111011010;assign rom[6609] = 'b111011010;assign rom[6610] = 'b111011010;assign rom[6611] = 'b111011000;assign rom[6612] = 'b111011000;assign rom[6613] = 'b111011000;assign rom[6614] = 'b111011000;assign rom[6615] = 'b101111000;assign rom[6616] = 'b000110011;assign rom[6617] = 'b110000010;assign rom[6618] = 'b001101010;assign rom[6619] = 'b001011000;assign rom[6620] = 'b101001000;assign rom[6621] = 'b000101011;assign rom[6622] = 'b110000010;assign rom[6623] = 'b111000000;assign rom[6624] = 'b101001100;assign rom[6625] = 'b001001010;assign rom[6626] = 'b111111000;assign rom[6627] = 'b111101000;assign rom[6628] = 'b101001111;assign rom[6629] = 'b000111010;assign rom[6630] = 'b101110110;assign rom[6631] = 'b101100010;assign rom[6632] = 'b101001100;assign rom[6633] = 'b001001010;assign rom[6634] = 'b111011010;assign rom[6635] = 'b111011010;assign rom[6636] = 'b111011010;assign rom[6637] = 'b111011010;assign rom[6638] = 'b111011000;assign rom[6639] = 'b111011000;assign rom[6640] = 'b111011000;assign rom[6641] = 'b111011000;assign rom[6642] = 'b101111000;assign rom[6643] = 'b000110011;assign rom[6644] = 'b110000010;assign rom[6645] = 'b001101010;assign rom[6646] = 'b001011000;assign rom[6647] = 'b101001000;assign rom[6648] = 'b000101011;assign rom[6649] = 'b110000010;assign rom[6650] = 'b111000000;assign rom[6651] = 'b101001100;assign rom[6652] = 'b001001010;assign rom[6653] = 'b111111000;assign rom[6654] = 'b111101000;assign rom[6655] = 'b101001111;assign rom[6656] = 'b000111010;assign rom[6657] = 'b101110110;assign rom[6658] = 'b101100010;assign rom[6659] = 'b101001100;assign rom[6660] = 'b001001010;assign rom[6661] = 'b111011010;assign rom[6662] = 'b111011010;assign rom[6663] = 'b111011010;assign rom[6664] = 'b111011010;assign rom[6665] = 'b111011000;assign rom[6666] = 'b111011000;assign rom[6667] = 'b111011000;assign rom[6668] = 'b111011000;assign rom[6669] = 'b101111000;assign rom[6670] = 'b000110011;assign rom[6671] = 'b110000010;assign rom[6672] = 'b001101010;assign rom[6673] = 'b001011000;assign rom[6674] = 'b101001000;assign rom[6675] = 'b000101011;assign rom[6676] = 'b110000010;assign rom[6677] = 'b111000000;assign rom[6678] = 'b101001100;assign rom[6679] = 'b001001010;assign rom[6680] = 'b111111000;assign rom[6681] = 'b111101000;assign rom[6682] = 'b101001111;assign rom[6683] = 'b000111010;assign rom[6684] = 'b101110110;assign rom[6685] = 'b101100010;assign rom[6686] = 'b101001100;assign rom[6687] = 'b001001010;assign rom[6688] = 'b111011010;assign rom[6689] = 'b111011010;assign rom[6690] = 'b111011010;assign rom[6691] = 'b111011010;assign rom[6692] = 'b111011000;assign rom[6693] = 'b111011000;assign rom[6694] = 'b111011000;assign rom[6695] = 'b111011000;assign rom[6696] = 'b101111000;assign rom[6697] = 'b000110011;assign rom[6698] = 'b110000010;assign rom[6699] = 'b001101010;assign rom[6700] = 'b001011000;assign rom[6701] = 'b101001000;assign rom[6702] = 'b000101011;assign rom[6703] = 'b110000010;assign rom[6704] = 'b111000000;assign rom[6705] = 'b101001100;assign rom[6706] = 'b001001010;assign rom[6707] = 'b111111000;assign rom[6708] = 'b111101000;assign rom[6709] = 'b101001111;assign rom[6710] = 'b000111010;assign rom[6711] = 'b101110110;assign rom[6712] = 'b101100010;assign rom[6713] = 'b101001100;assign rom[6714] = 'b001001010;assign rom[6715] = 'b111011010;assign rom[6716] = 'b111011010;assign rom[6717] = 'b111011010;assign rom[6718] = 'b111011010;assign rom[6719] = 'b111011000;assign rom[6720] = 'b111011000;assign rom[6721] = 'b111011000;assign rom[6722] = 'b111011000;assign rom[6723] = 'b101111000;assign rom[6724] = 'b000110011;assign rom[6725] = 'b110000010;assign rom[6726] = 'b001101010;assign rom[6727] = 'b001011000;assign rom[6728] = 'b101001000;assign rom[6729] = 'b000101011;assign rom[6730] = 'b110000010;assign rom[6731] = 'b111000000;assign rom[6732] = 'b101001100;assign rom[6733] = 'b001001010;assign rom[6734] = 'b111111000;assign rom[6735] = 'b111101000;assign rom[6736] = 'b101001111;assign rom[6737] = 'b000111010;assign rom[6738] = 'b101110110;assign rom[6739] = 'b101100010;assign rom[6740] = 'b101001100;assign rom[6741] = 'b001001010;assign rom[6742] = 'b111011010;assign rom[6743] = 'b111011010;assign rom[6744] = 'b111011010;assign rom[6745] = 'b111011010;assign rom[6746] = 'b111011000;assign rom[6747] = 'b111011000;assign rom[6748] = 'b111011000;assign rom[6749] = 'b111011000;assign rom[6750] = 'b101111000;assign rom[6751] = 'b000110011;assign rom[6752] = 'b110000010;assign rom[6753] = 'b001101010;assign rom[6754] = 'b001011000;assign rom[6755] = 'b101001000;assign rom[6756] = 'b000101011;assign rom[6757] = 'b110000010;assign rom[6758] = 'b111000000;assign rom[6759] = 'b101001100;assign rom[6760] = 'b001001010;assign rom[6761] = 'b001000110;assign rom[6762] = 'b001100100;assign rom[6763] = 'b101100010;assign rom[6764] = 'b101001100;assign rom[6765] = 'b001001010;assign rom[6766] = 'b111011010;assign rom[6767] = 'b111011010;assign rom[6768] = 'b111011010;assign rom[6769] = 'b111011010;assign rom[6770] = 'b111011000;assign rom[6771] = 'b111011000;assign rom[6772] = 'b111011000;assign rom[6773] = 'b111011000;assign rom[6774] = 'b101111000;assign rom[6775] = 'b000110011;assign rom[6776] = 'b110000010;assign rom[6777] = 'b001101010;assign rom[6778] = 'b001011000;assign rom[6779] = 'b101001000;assign rom[6780] = 'b000101011;assign rom[6781] = 'b110000010;assign rom[6782] = 'b111000000;assign rom[6783] = 'b101001100;assign rom[6784] = 'b001001010;assign rom[6785] = 'b111111000;assign rom[6786] = 'b111101000;assign rom[6787] = 'b101001111;assign rom[6788] = 'b000111010;assign rom[6789] = 'b101110110;assign rom[6790] = 'b101100010;assign rom[6791] = 'b101001100;assign rom[6792] = 'b001001010;assign rom[6793] = 'b111011010;assign rom[6794] = 'b111011010;assign rom[6795] = 'b111011010;assign rom[6796] = 'b111011010;assign rom[6797] = 'b111011000;assign rom[6798] = 'b111011000;assign rom[6799] = 'b111011000;assign rom[6800] = 'b111011000;assign rom[6801] = 'b101111000;assign rom[6802] = 'b000110011;assign rom[6803] = 'b110000010;assign rom[6804] = 'b001101010;assign rom[6805] = 'b001011000;assign rom[6806] = 'b101001000;assign rom[6807] = 'b000101011;assign rom[6808] = 'b110000010;assign rom[6809] = 'b111000000;assign rom[6810] = 'b101001100;assign rom[6811] = 'b001001010;assign rom[6812] = 'b111111000;assign rom[6813] = 'b111101000;assign rom[6814] = 'b101001111;assign rom[6815] = 'b000111010;assign rom[6816] = 'b101110110;assign rom[6817] = 'b101100010;assign rom[6818] = 'b101001100;assign rom[6819] = 'b001001010;assign rom[6820] = 'b111011010;assign rom[6821] = 'b111011010;assign rom[6822] = 'b111011010;assign rom[6823] = 'b111011010;assign rom[6824] = 'b111011000;assign rom[6825] = 'b111011000;assign rom[6826] = 'b111011000;assign rom[6827] = 'b111011000;assign rom[6828] = 'b101111000;assign rom[6829] = 'b000110011;assign rom[6830] = 'b110000010;assign rom[6831] = 'b001101010;assign rom[6832] = 'b001011000;assign rom[6833] = 'b101001000;assign rom[6834] = 'b000101011;assign rom[6835] = 'b110000010;assign rom[6836] = 'b111000000;assign rom[6837] = 'b101001100;assign rom[6838] = 'b001001010;assign rom[6839] = 'b111111000;assign rom[6840] = 'b111101000;assign rom[6841] = 'b101001111;assign rom[6842] = 'b000111010;assign rom[6843] = 'b101110110;assign rom[6844] = 'b101100010;assign rom[6845] = 'b101001100;assign rom[6846] = 'b001001010;assign rom[6847] = 'b111011010;assign rom[6848] = 'b111011010;assign rom[6849] = 'b111011010;assign rom[6850] = 'b111011010;assign rom[6851] = 'b111011000;assign rom[6852] = 'b111011000;assign rom[6853] = 'b111011000;assign rom[6854] = 'b111011000;assign rom[6855] = 'b101111000;assign rom[6856] = 'b000110011;assign rom[6857] = 'b110000010;assign rom[6858] = 'b001101010;assign rom[6859] = 'b001011000;assign rom[6860] = 'b101001000;assign rom[6861] = 'b000101011;assign rom[6862] = 'b110000010;assign rom[6863] = 'b111000000;assign rom[6864] = 'b101001100;assign rom[6865] = 'b001001010;assign rom[6866] = 'b111111000;assign rom[6867] = 'b111101000;assign rom[6868] = 'b101001111;assign rom[6869] = 'b000111010;assign rom[6870] = 'b101110110;assign rom[6871] = 'b101100010;assign rom[6872] = 'b101001100;assign rom[6873] = 'b001001010;assign rom[6874] = 'b111011010;assign rom[6875] = 'b111011010;assign rom[6876] = 'b111011010;assign rom[6877] = 'b111011010;assign rom[6878] = 'b111011000;assign rom[6879] = 'b111011000;assign rom[6880] = 'b111011000;assign rom[6881] = 'b111011000;assign rom[6882] = 'b101111000;assign rom[6883] = 'b000110011;assign rom[6884] = 'b110000010;assign rom[6885] = 'b001101010;assign rom[6886] = 'b001011000;assign rom[6887] = 'b101001000;assign rom[6888] = 'b000101011;assign rom[6889] = 'b110000010;assign rom[6890] = 'b111000000;assign rom[6891] = 'b101001100;assign rom[6892] = 'b001001010;assign rom[6893] = 'b111111000;assign rom[6894] = 'b111101000;assign rom[6895] = 'b101001111;assign rom[6896] = 'b000111010;assign rom[6897] = 'b101110110;assign rom[6898] = 'b101100010;assign rom[6899] = 'b101001100;assign rom[6900] = 'b001001010;assign rom[6901] = 'b111011010;assign rom[6902] = 'b111011010;assign rom[6903] = 'b111011010;assign rom[6904] = 'b111011010;assign rom[6905] = 'b111011000;assign rom[6906] = 'b111011000;assign rom[6907] = 'b111011000;assign rom[6908] = 'b111011000;assign rom[6909] = 'b101111000;assign rom[6910] = 'b000110011;assign rom[6911] = 'b110000010;assign rom[6912] = 'b001101010;assign rom[6913] = 'b001011000;assign rom[6914] = 'b101001000;assign rom[6915] = 'b000101011;assign rom[6916] = 'b110000010;assign rom[6917] = 'b111000000;assign rom[6918] = 'b101001100;assign rom[6919] = 'b001001010;assign rom[6920] = 'b111111000;assign rom[6921] = 'b111101000;assign rom[6922] = 'b101001111;assign rom[6923] = 'b000111010;assign rom[6924] = 'b101110110;assign rom[6925] = 'b101100010;assign rom[6926] = 'b101001100;assign rom[6927] = 'b001001010;assign rom[6928] = 'b111011010;assign rom[6929] = 'b111011010;assign rom[6930] = 'b111011010;assign rom[6931] = 'b111011010;assign rom[6932] = 'b111011000;assign rom[6933] = 'b111011000;assign rom[6934] = 'b111011000;assign rom[6935] = 'b111011000;assign rom[6936] = 'b101111000;assign rom[6937] = 'b000110011;assign rom[6938] = 'b110000010;assign rom[6939] = 'b001101010;assign rom[6940] = 'b001011000;assign rom[6941] = 'b101001000;assign rom[6942] = 'b000101011;assign rom[6943] = 'b110000010;assign rom[6944] = 'b111000000;assign rom[6945] = 'b101001100;assign rom[6946] = 'b001001010;assign rom[6947] = 'b111111000;assign rom[6948] = 'b111101000;assign rom[6949] = 'b101001111;assign rom[6950] = 'b000111010;assign rom[6951] = 'b101110110;assign rom[6952] = 'b101100010;assign rom[6953] = 'b101001100;assign rom[6954] = 'b001001010;assign rom[6955] = 'b111011010;assign rom[6956] = 'b111011010;assign rom[6957] = 'b111011010;assign rom[6958] = 'b111011010;assign rom[6959] = 'b111011000;assign rom[6960] = 'b111011000;assign rom[6961] = 'b111011000;assign rom[6962] = 'b111011000;assign rom[6963] = 'b101111000;assign rom[6964] = 'b000110011;assign rom[6965] = 'b110000010;assign rom[6966] = 'b001101010;assign rom[6967] = 'b001011000;assign rom[6968] = 'b101001000;assign rom[6969] = 'b000101011;assign rom[6970] = 'b110000010;assign rom[6971] = 'b111000000;assign rom[6972] = 'b101001100;assign rom[6973] = 'b001001010;assign rom[6974] = 'b111111000;assign rom[6975] = 'b111101000;assign rom[6976] = 'b101001111;assign rom[6977] = 'b000111010;assign rom[6978] = 'b101110110;assign rom[6979] = 'b101100010;assign rom[6980] = 'b101001100;assign rom[6981] = 'b001001010;assign rom[6982] = 'b111011010;assign rom[6983] = 'b111011010;assign rom[6984] = 'b111011010;assign rom[6985] = 'b111011010;assign rom[6986] = 'b111011000;assign rom[6987] = 'b111011000;assign rom[6988] = 'b111011000;assign rom[6989] = 'b111011000;assign rom[6990] = 'b101111000;assign rom[6991] = 'b000110011;assign rom[6992] = 'b110000010;assign rom[6993] = 'b001101010;assign rom[6994] = 'b001011000;assign rom[6995] = 'b101001000;assign rom[6996] = 'b000101011;assign rom[6997] = 'b110000010;assign rom[6998] = 'b111000000;assign rom[6999] = 'b101001100;assign rom[7000] = 'b001001010;assign rom[7001] = 'b001000110;assign rom[7002] = 'b001100100;assign rom[7003] = 'b101100010;assign rom[7004] = 'b101001100;assign rom[7005] = 'b001001010;assign rom[7006] = 'b111011010;assign rom[7007] = 'b111011010;assign rom[7008] = 'b111011010;assign rom[7009] = 'b111011010;assign rom[7010] = 'b111011000;assign rom[7011] = 'b111011000;assign rom[7012] = 'b111011000;assign rom[7013] = 'b111011000;assign rom[7014] = 'b101111000;assign rom[7015] = 'b000110011;assign rom[7016] = 'b110000010;assign rom[7017] = 'b001101010;assign rom[7018] = 'b001011000;assign rom[7019] = 'b101001000;assign rom[7020] = 'b000101011;assign rom[7021] = 'b110000010;assign rom[7022] = 'b111000000;assign rom[7023] = 'b101001100;assign rom[7024] = 'b001001010;assign rom[7025] = 'b111111000;assign rom[7026] = 'b111101000;assign rom[7027] = 'b101001111;assign rom[7028] = 'b000111010;assign rom[7029] = 'b101110110;assign rom[7030] = 'b101100010;assign rom[7031] = 'b101001100;assign rom[7032] = 'b001001010;assign rom[7033] = 'b111011010;assign rom[7034] = 'b111011010;assign rom[7035] = 'b111011010;assign rom[7036] = 'b111011010;assign rom[7037] = 'b111011000;assign rom[7038] = 'b111011000;assign rom[7039] = 'b111011000;assign rom[7040] = 'b111011000;assign rom[7041] = 'b101111000;assign rom[7042] = 'b000110011;assign rom[7043] = 'b110000010;assign rom[7044] = 'b001101010;assign rom[7045] = 'b001011000;assign rom[7046] = 'b101001000;assign rom[7047] = 'b000101011;assign rom[7048] = 'b110000010;assign rom[7049] = 'b111000000;assign rom[7050] = 'b101001100;assign rom[7051] = 'b001001010;assign rom[7052] = 'b111111000;assign rom[7053] = 'b111101000;assign rom[7054] = 'b101001111;assign rom[7055] = 'b000111010;assign rom[7056] = 'b101110110;assign rom[7057] = 'b101100010;assign rom[7058] = 'b101001100;assign rom[7059] = 'b001001010;assign rom[7060] = 'b111011010;assign rom[7061] = 'b111011010;assign rom[7062] = 'b111011010;assign rom[7063] = 'b111011010;assign rom[7064] = 'b111011000;assign rom[7065] = 'b111011000;assign rom[7066] = 'b111011000;assign rom[7067] = 'b111011000;assign rom[7068] = 'b101111000;assign rom[7069] = 'b000110011;assign rom[7070] = 'b110000010;assign rom[7071] = 'b001101010;assign rom[7072] = 'b001011000;assign rom[7073] = 'b101001000;assign rom[7074] = 'b000101011;assign rom[7075] = 'b110000010;assign rom[7076] = 'b111000000;assign rom[7077] = 'b101001100;assign rom[7078] = 'b001001010;assign rom[7079] = 'b111111000;assign rom[7080] = 'b111101000;assign rom[7081] = 'b101001111;assign rom[7082] = 'b000111010;assign rom[7083] = 'b101110110;assign rom[7084] = 'b101100010;assign rom[7085] = 'b101001100;assign rom[7086] = 'b001001010;assign rom[7087] = 'b111011010;assign rom[7088] = 'b111011010;assign rom[7089] = 'b111011010;assign rom[7090] = 'b111011010;assign rom[7091] = 'b111011000;assign rom[7092] = 'b111011000;assign rom[7093] = 'b111011000;assign rom[7094] = 'b111011000;assign rom[7095] = 'b101111000;assign rom[7096] = 'b000110011;assign rom[7097] = 'b110000010;assign rom[7098] = 'b001101010;assign rom[7099] = 'b001011000;assign rom[7100] = 'b101001000;assign rom[7101] = 'b000101011;assign rom[7102] = 'b110000010;assign rom[7103] = 'b111000000;assign rom[7104] = 'b101001100;assign rom[7105] = 'b001001010;assign rom[7106] = 'b111111000;assign rom[7107] = 'b111101000;assign rom[7108] = 'b101001111;assign rom[7109] = 'b000111010;assign rom[7110] = 'b101110110;assign rom[7111] = 'b101100010;assign rom[7112] = 'b101001100;assign rom[7113] = 'b001001010;assign rom[7114] = 'b111011010;assign rom[7115] = 'b111011010;assign rom[7116] = 'b111011010;assign rom[7117] = 'b111011010;assign rom[7118] = 'b111011000;assign rom[7119] = 'b111011000;assign rom[7120] = 'b111011000;assign rom[7121] = 'b111011000;assign rom[7122] = 'b101111000;assign rom[7123] = 'b000110011;assign rom[7124] = 'b110000010;assign rom[7125] = 'b001101010;assign rom[7126] = 'b001011000;assign rom[7127] = 'b101001000;assign rom[7128] = 'b000101011;assign rom[7129] = 'b110000010;assign rom[7130] = 'b111000000;assign rom[7131] = 'b101001100;assign rom[7132] = 'b001001010;assign rom[7133] = 'b111111000;assign rom[7134] = 'b111101000;assign rom[7135] = 'b101001111;assign rom[7136] = 'b000111010;assign rom[7137] = 'b101110110;assign rom[7138] = 'b101100010;assign rom[7139] = 'b101001100;assign rom[7140] = 'b001001010;assign rom[7141] = 'b111011010;assign rom[7142] = 'b111011010;assign rom[7143] = 'b111011010;assign rom[7144] = 'b111011010;assign rom[7145] = 'b111011000;assign rom[7146] = 'b111011000;assign rom[7147] = 'b111011000;assign rom[7148] = 'b111011000;assign rom[7149] = 'b101111000;assign rom[7150] = 'b000110011;assign rom[7151] = 'b110000010;assign rom[7152] = 'b001101010;assign rom[7153] = 'b001011000;assign rom[7154] = 'b101001000;assign rom[7155] = 'b000101011;assign rom[7156] = 'b110000010;assign rom[7157] = 'b111000000;assign rom[7158] = 'b101001100;assign rom[7159] = 'b001001010;assign rom[7160] = 'b111111000;assign rom[7161] = 'b111101000;assign rom[7162] = 'b101001111;assign rom[7163] = 'b000111010;assign rom[7164] = 'b101110110;assign rom[7165] = 'b101100010;assign rom[7166] = 'b101001100;assign rom[7167] = 'b001001010;assign rom[7168] = 'b111011010;assign rom[7169] = 'b111011010;assign rom[7170] = 'b111011010;assign rom[7171] = 'b111011010;assign rom[7172] = 'b111011000;assign rom[7173] = 'b111011000;assign rom[7174] = 'b111011000;assign rom[7175] = 'b111011000;assign rom[7176] = 'b101111000;assign rom[7177] = 'b000110011;assign rom[7178] = 'b110000010;assign rom[7179] = 'b001101010;assign rom[7180] = 'b001011000;assign rom[7181] = 'b101001000;assign rom[7182] = 'b000101011;assign rom[7183] = 'b110000010;assign rom[7184] = 'b111000000;assign rom[7185] = 'b101001100;assign rom[7186] = 'b001001010;assign rom[7187] = 'b111111000;assign rom[7188] = 'b111101000;assign rom[7189] = 'b101001111;assign rom[7190] = 'b000111010;assign rom[7191] = 'b101110110;assign rom[7192] = 'b101100010;assign rom[7193] = 'b101001100;assign rom[7194] = 'b001001010;assign rom[7195] = 'b111011010;assign rom[7196] = 'b111011010;assign rom[7197] = 'b111011010;assign rom[7198] = 'b111011010;assign rom[7199] = 'b111011000;assign rom[7200] = 'b111011000;assign rom[7201] = 'b111011000;assign rom[7202] = 'b111011000;assign rom[7203] = 'b101111000;assign rom[7204] = 'b000110011;assign rom[7205] = 'b110000010;assign rom[7206] = 'b001101010;assign rom[7207] = 'b001011000;assign rom[7208] = 'b101001000;assign rom[7209] = 'b000101011;assign rom[7210] = 'b110000010;assign rom[7211] = 'b111000000;assign rom[7212] = 'b101001100;assign rom[7213] = 'b001001010;assign rom[7214] = 'b111111000;assign rom[7215] = 'b111101000;assign rom[7216] = 'b101001111;assign rom[7217] = 'b000111010;assign rom[7218] = 'b101110110;assign rom[7219] = 'b101100010;assign rom[7220] = 'b101001100;assign rom[7221] = 'b001001010;assign rom[7222] = 'b111011010;assign rom[7223] = 'b111011010;assign rom[7224] = 'b111011010;assign rom[7225] = 'b111011010;assign rom[7226] = 'b111011000;assign rom[7227] = 'b111011000;assign rom[7228] = 'b111011000;assign rom[7229] = 'b111011000;assign rom[7230] = 'b101111000;assign rom[7231] = 'b000110011;assign rom[7232] = 'b110000010;assign rom[7233] = 'b001101010;assign rom[7234] = 'b001011000;assign rom[7235] = 'b101001000;assign rom[7236] = 'b000101011;assign rom[7237] = 'b110000010;assign rom[7238] = 'b111000000;assign rom[7239] = 'b101001100;assign rom[7240] = 'b001001010;assign rom[7241] = 'b001000110;assign rom[7242] = 'b001100100;assign rom[7243] = 'b101100010;assign rom[7244] = 'b101001100;assign rom[7245] = 'b001001010;assign rom[7246] = 'b111011010;assign rom[7247] = 'b111011010;assign rom[7248] = 'b111011010;assign rom[7249] = 'b111011010;assign rom[7250] = 'b111011000;assign rom[7251] = 'b111011000;assign rom[7252] = 'b111011000;assign rom[7253] = 'b111011000;assign rom[7254] = 'b101111000;assign rom[7255] = 'b000110011;assign rom[7256] = 'b110000010;assign rom[7257] = 'b001101010;assign rom[7258] = 'b001011000;assign rom[7259] = 'b101001000;assign rom[7260] = 'b000101011;assign rom[7261] = 'b110000010;assign rom[7262] = 'b111000000;assign rom[7263] = 'b101001100;assign rom[7264] = 'b001001010;assign rom[7265] = 'b111111000;assign rom[7266] = 'b111101000;assign rom[7267] = 'b101001111;assign rom[7268] = 'b000111010;assign rom[7269] = 'b101110110;assign rom[7270] = 'b101100010;assign rom[7271] = 'b101001100;assign rom[7272] = 'b001001010;assign rom[7273] = 'b111011010;assign rom[7274] = 'b111011010;assign rom[7275] = 'b111011010;assign rom[7276] = 'b111011010;assign rom[7277] = 'b111011000;assign rom[7278] = 'b111011000;assign rom[7279] = 'b111011000;assign rom[7280] = 'b111011000;assign rom[7281] = 'b101111000;assign rom[7282] = 'b000110011;assign rom[7283] = 'b110000010;assign rom[7284] = 'b001101010;assign rom[7285] = 'b001011000;assign rom[7286] = 'b101001000;assign rom[7287] = 'b000101011;assign rom[7288] = 'b110000010;assign rom[7289] = 'b111000000;assign rom[7290] = 'b101001100;assign rom[7291] = 'b001001010;assign rom[7292] = 'b111111000;assign rom[7293] = 'b111101000;assign rom[7294] = 'b101001111;assign rom[7295] = 'b000111010;assign rom[7296] = 'b101110110;assign rom[7297] = 'b101100010;assign rom[7298] = 'b101001100;assign rom[7299] = 'b001001010;assign rom[7300] = 'b111011010;assign rom[7301] = 'b111011010;assign rom[7302] = 'b111011010;assign rom[7303] = 'b111011010;assign rom[7304] = 'b111011000;assign rom[7305] = 'b111011000;assign rom[7306] = 'b111011000;assign rom[7307] = 'b111011000;assign rom[7308] = 'b101111000;assign rom[7309] = 'b000110011;assign rom[7310] = 'b110000010;assign rom[7311] = 'b001101010;assign rom[7312] = 'b001011000;assign rom[7313] = 'b101001000;assign rom[7314] = 'b000101011;assign rom[7315] = 'b110000010;assign rom[7316] = 'b111000000;assign rom[7317] = 'b101001100;assign rom[7318] = 'b001001010;assign rom[7319] = 'b111111000;assign rom[7320] = 'b111101000;assign rom[7321] = 'b101001111;assign rom[7322] = 'b000111010;assign rom[7323] = 'b101110110;assign rom[7324] = 'b101100010;assign rom[7325] = 'b101001100;assign rom[7326] = 'b001001010;assign rom[7327] = 'b111011010;assign rom[7328] = 'b111011010;assign rom[7329] = 'b111011010;assign rom[7330] = 'b111011010;assign rom[7331] = 'b111011000;assign rom[7332] = 'b111011000;assign rom[7333] = 'b111011000;assign rom[7334] = 'b111011000;assign rom[7335] = 'b101111000;assign rom[7336] = 'b000110011;assign rom[7337] = 'b110000010;assign rom[7338] = 'b001101010;assign rom[7339] = 'b001011000;assign rom[7340] = 'b101001000;assign rom[7341] = 'b000101011;assign rom[7342] = 'b110000010;assign rom[7343] = 'b111000000;assign rom[7344] = 'b101001100;assign rom[7345] = 'b001001010;assign rom[7346] = 'b111111000;assign rom[7347] = 'b111101000;assign rom[7348] = 'b101001111;assign rom[7349] = 'b000111010;assign rom[7350] = 'b101110110;assign rom[7351] = 'b101100010;assign rom[7352] = 'b101001100;assign rom[7353] = 'b001001010;assign rom[7354] = 'b111011010;assign rom[7355] = 'b111011010;assign rom[7356] = 'b111011010;assign rom[7357] = 'b111011010;assign rom[7358] = 'b111011000;assign rom[7359] = 'b111011000;assign rom[7360] = 'b111011000;assign rom[7361] = 'b111011000;assign rom[7362] = 'b101111000;assign rom[7363] = 'b000110011;assign rom[7364] = 'b110000010;assign rom[7365] = 'b001101010;assign rom[7366] = 'b001011000;assign rom[7367] = 'b101001000;assign rom[7368] = 'b000101011;assign rom[7369] = 'b110000010;assign rom[7370] = 'b111000000;assign rom[7371] = 'b101001100;assign rom[7372] = 'b001001010;assign rom[7373] = 'b111111000;assign rom[7374] = 'b111101000;assign rom[7375] = 'b101001111;assign rom[7376] = 'b000111010;assign rom[7377] = 'b101110110;assign rom[7378] = 'b101100010;assign rom[7379] = 'b101001100;assign rom[7380] = 'b001001010;assign rom[7381] = 'b111011010;assign rom[7382] = 'b111011010;assign rom[7383] = 'b111011010;assign rom[7384] = 'b111011010;assign rom[7385] = 'b111011000;assign rom[7386] = 'b111011000;assign rom[7387] = 'b111011000;assign rom[7388] = 'b111011000;assign rom[7389] = 'b101111000;assign rom[7390] = 'b000110011;assign rom[7391] = 'b110000010;assign rom[7392] = 'b001101010;assign rom[7393] = 'b001011000;assign rom[7394] = 'b101001000;assign rom[7395] = 'b000101011;assign rom[7396] = 'b110000010;assign rom[7397] = 'b111000000;assign rom[7398] = 'b101001100;assign rom[7399] = 'b001001010;assign rom[7400] = 'b111111000;assign rom[7401] = 'b111101000;assign rom[7402] = 'b101001111;assign rom[7403] = 'b000111010;assign rom[7404] = 'b101110110;assign rom[7405] = 'b101100010;assign rom[7406] = 'b101001100;assign rom[7407] = 'b001001010;assign rom[7408] = 'b111011010;assign rom[7409] = 'b111011010;assign rom[7410] = 'b111011010;assign rom[7411] = 'b111011010;assign rom[7412] = 'b111011000;assign rom[7413] = 'b111011000;assign rom[7414] = 'b111011000;assign rom[7415] = 'b111011000;assign rom[7416] = 'b101111000;assign rom[7417] = 'b000110011;assign rom[7418] = 'b110000010;assign rom[7419] = 'b001101010;assign rom[7420] = 'b001011000;assign rom[7421] = 'b101001000;assign rom[7422] = 'b000101011;assign rom[7423] = 'b110000010;assign rom[7424] = 'b111000000;assign rom[7425] = 'b101001100;assign rom[7426] = 'b001001010;assign rom[7427] = 'b111111000;assign rom[7428] = 'b111101000;assign rom[7429] = 'b101001111;assign rom[7430] = 'b000111010;assign rom[7431] = 'b101110110;assign rom[7432] = 'b101100010;assign rom[7433] = 'b101001100;assign rom[7434] = 'b001001010;assign rom[7435] = 'b111011010;assign rom[7436] = 'b111011010;assign rom[7437] = 'b111011010;assign rom[7438] = 'b111011010;assign rom[7439] = 'b111011000;assign rom[7440] = 'b111011000;assign rom[7441] = 'b111011000;assign rom[7442] = 'b111011000;assign rom[7443] = 'b101111000;assign rom[7444] = 'b000110011;assign rom[7445] = 'b110000010;assign rom[7446] = 'b001101010;assign rom[7447] = 'b001011000;assign rom[7448] = 'b101001000;assign rom[7449] = 'b000101011;assign rom[7450] = 'b110000010;assign rom[7451] = 'b111000000;assign rom[7452] = 'b101001100;assign rom[7453] = 'b001001010;assign rom[7454] = 'b111111000;assign rom[7455] = 'b111101000;assign rom[7456] = 'b101001111;assign rom[7457] = 'b000111010;assign rom[7458] = 'b101110110;assign rom[7459] = 'b101100010;assign rom[7460] = 'b101001100;assign rom[7461] = 'b001001010;assign rom[7462] = 'b111011010;assign rom[7463] = 'b111011010;assign rom[7464] = 'b111011010;assign rom[7465] = 'b111011010;assign rom[7466] = 'b111011000;assign rom[7467] = 'b111011000;assign rom[7468] = 'b111011000;assign rom[7469] = 'b111011000;assign rom[7470] = 'b101111000;assign rom[7471] = 'b000110011;assign rom[7472] = 'b110000010;assign rom[7473] = 'b001101010;assign rom[7474] = 'b001011000;assign rom[7475] = 'b101001000;assign rom[7476] = 'b000101011;assign rom[7477] = 'b110000010;assign rom[7478] = 'b111000000;assign rom[7479] = 'b101001100;assign rom[7480] = 'b001001010;assign rom[7481] = 'b001000110;assign rom[7482] = 'b001100100;assign rom[7483] = 'b101100010;assign rom[7484] = 'b101001100;assign rom[7485] = 'b001001010;assign rom[7486] = 'b111011010;assign rom[7487] = 'b111011010;assign rom[7488] = 'b111011010;assign rom[7489] = 'b111011010;assign rom[7490] = 'b111011000;assign rom[7491] = 'b111011000;assign rom[7492] = 'b111011000;assign rom[7493] = 'b111011000;assign rom[7494] = 'b101111000;assign rom[7495] = 'b000110011;assign rom[7496] = 'b110000010;assign rom[7497] = 'b001101010;assign rom[7498] = 'b001011000;assign rom[7499] = 'b101001000;assign rom[7500] = 'b000101011;assign rom[7501] = 'b110000010;assign rom[7502] = 'b111000000;assign rom[7503] = 'b101001100;assign rom[7504] = 'b001001010;assign rom[7505] = 'b111111000;assign rom[7506] = 'b111101000;assign rom[7507] = 'b101001111;assign rom[7508] = 'b000111010;assign rom[7509] = 'b101110110;assign rom[7510] = 'b101100010;assign rom[7511] = 'b101001100;assign rom[7512] = 'b001001010;assign rom[7513] = 'b111011010;assign rom[7514] = 'b111011010;assign rom[7515] = 'b111011010;assign rom[7516] = 'b111011010;assign rom[7517] = 'b111011000;assign rom[7518] = 'b111011000;assign rom[7519] = 'b111011000;assign rom[7520] = 'b111011000;assign rom[7521] = 'b101111000;assign rom[7522] = 'b000110011;assign rom[7523] = 'b110000010;assign rom[7524] = 'b001101010;assign rom[7525] = 'b001011000;assign rom[7526] = 'b101001000;assign rom[7527] = 'b000101011;assign rom[7528] = 'b110000010;assign rom[7529] = 'b111000000;assign rom[7530] = 'b101001100;assign rom[7531] = 'b001001010;assign rom[7532] = 'b111111000;assign rom[7533] = 'b111101000;assign rom[7534] = 'b101001111;assign rom[7535] = 'b000111010;assign rom[7536] = 'b101110110;assign rom[7537] = 'b101100010;assign rom[7538] = 'b101001100;assign rom[7539] = 'b001001010;assign rom[7540] = 'b111011010;assign rom[7541] = 'b111011010;assign rom[7542] = 'b111011010;assign rom[7543] = 'b111011010;assign rom[7544] = 'b111011000;assign rom[7545] = 'b111011000;assign rom[7546] = 'b111011000;assign rom[7547] = 'b111011000;assign rom[7548] = 'b101111000;assign rom[7549] = 'b000110011;assign rom[7550] = 'b110000010;assign rom[7551] = 'b001101010;assign rom[7552] = 'b001011000;assign rom[7553] = 'b101001000;assign rom[7554] = 'b000101011;assign rom[7555] = 'b110000010;assign rom[7556] = 'b111000000;assign rom[7557] = 'b101001100;assign rom[7558] = 'b001001010;assign rom[7559] = 'b111111000;assign rom[7560] = 'b111101000;assign rom[7561] = 'b101001111;assign rom[7562] = 'b000111010;assign rom[7563] = 'b101110110;assign rom[7564] = 'b101100010;assign rom[7565] = 'b101001100;assign rom[7566] = 'b001001010;assign rom[7567] = 'b111011010;assign rom[7568] = 'b111011010;assign rom[7569] = 'b111011010;assign rom[7570] = 'b111011010;assign rom[7571] = 'b111011000;assign rom[7572] = 'b111011000;assign rom[7573] = 'b111011000;assign rom[7574] = 'b111011000;assign rom[7575] = 'b101111000;assign rom[7576] = 'b000110011;assign rom[7577] = 'b110000010;assign rom[7578] = 'b001101010;assign rom[7579] = 'b001011000;assign rom[7580] = 'b101001000;assign rom[7581] = 'b000101011;assign rom[7582] = 'b110000010;assign rom[7583] = 'b111000000;assign rom[7584] = 'b101001100;assign rom[7585] = 'b001001010;assign rom[7586] = 'b111111000;assign rom[7587] = 'b111101000;assign rom[7588] = 'b101001111;assign rom[7589] = 'b000111010;assign rom[7590] = 'b101110110;assign rom[7591] = 'b101100010;assign rom[7592] = 'b101001100;assign rom[7593] = 'b001001010;assign rom[7594] = 'b111011010;assign rom[7595] = 'b111011010;assign rom[7596] = 'b111011010;assign rom[7597] = 'b111011010;assign rom[7598] = 'b111011000;assign rom[7599] = 'b111011000;assign rom[7600] = 'b111011000;assign rom[7601] = 'b111011000;assign rom[7602] = 'b101111000;assign rom[7603] = 'b000110011;assign rom[7604] = 'b110000010;assign rom[7605] = 'b001101010;assign rom[7606] = 'b001011000;assign rom[7607] = 'b101001000;assign rom[7608] = 'b000101011;assign rom[7609] = 'b110000010;assign rom[7610] = 'b111000000;assign rom[7611] = 'b101001100;assign rom[7612] = 'b001001010;assign rom[7613] = 'b111111000;assign rom[7614] = 'b111101000;assign rom[7615] = 'b101001111;assign rom[7616] = 'b000111010;assign rom[7617] = 'b101110110;assign rom[7618] = 'b101100010;assign rom[7619] = 'b101001100;assign rom[7620] = 'b001001010;assign rom[7621] = 'b111011010;assign rom[7622] = 'b111011010;assign rom[7623] = 'b111011010;assign rom[7624] = 'b111011010;assign rom[7625] = 'b111011000;assign rom[7626] = 'b111011000;assign rom[7627] = 'b111011000;assign rom[7628] = 'b111011000;assign rom[7629] = 'b101111000;assign rom[7630] = 'b000110011;assign rom[7631] = 'b110000010;assign rom[7632] = 'b001101010;assign rom[7633] = 'b001011000;assign rom[7634] = 'b101001000;assign rom[7635] = 'b000101011;assign rom[7636] = 'b110000010;assign rom[7637] = 'b111000000;assign rom[7638] = 'b101001100;assign rom[7639] = 'b001001010;assign rom[7640] = 'b111111000;assign rom[7641] = 'b111101000;assign rom[7642] = 'b101001111;assign rom[7643] = 'b000111010;assign rom[7644] = 'b101110110;assign rom[7645] = 'b101100010;assign rom[7646] = 'b101001100;assign rom[7647] = 'b001001010;assign rom[7648] = 'b111011010;assign rom[7649] = 'b111011010;assign rom[7650] = 'b111011010;assign rom[7651] = 'b111011010;assign rom[7652] = 'b111011000;assign rom[7653] = 'b111011000;assign rom[7654] = 'b111011000;assign rom[7655] = 'b111011000;assign rom[7656] = 'b101111000;assign rom[7657] = 'b000110011;assign rom[7658] = 'b110000010;assign rom[7659] = 'b001101010;assign rom[7660] = 'b001011000;assign rom[7661] = 'b101001000;assign rom[7662] = 'b000101011;assign rom[7663] = 'b110000010;assign rom[7664] = 'b111000000;assign rom[7665] = 'b101001100;assign rom[7666] = 'b001001010;assign rom[7667] = 'b111111000;assign rom[7668] = 'b111101000;assign rom[7669] = 'b101001111;assign rom[7670] = 'b000111010;assign rom[7671] = 'b101110110;assign rom[7672] = 'b101100010;assign rom[7673] = 'b101001100;assign rom[7674] = 'b001001010;assign rom[7675] = 'b111011010;assign rom[7676] = 'b111011010;assign rom[7677] = 'b111011010;assign rom[7678] = 'b111011010;assign rom[7679] = 'b111011000;assign rom[7680] = 'b111011000;assign rom[7681] = 'b111011000;assign rom[7682] = 'b111011000;assign rom[7683] = 'b101111000;assign rom[7684] = 'b000110011;assign rom[7685] = 'b110000010;assign rom[7686] = 'b001101010;assign rom[7687] = 'b001011000;assign rom[7688] = 'b101001000;assign rom[7689] = 'b000101011;assign rom[7690] = 'b110000010;assign rom[7691] = 'b111000000;assign rom[7692] = 'b101001100;assign rom[7693] = 'b001001010;assign rom[7694] = 'b111111000;assign rom[7695] = 'b111101000;assign rom[7696] = 'b101001111;assign rom[7697] = 'b000111010;assign rom[7698] = 'b101110110;assign rom[7699] = 'b101100010;assign rom[7700] = 'b101001100;assign rom[7701] = 'b001001010;assign rom[7702] = 'b111011010;assign rom[7703] = 'b111011010;assign rom[7704] = 'b111011010;assign rom[7705] = 'b111011010;assign rom[7706] = 'b111011000;assign rom[7707] = 'b111011000;assign rom[7708] = 'b111011000;assign rom[7709] = 'b111011000;assign rom[7710] = 'b101111000;assign rom[7711] = 'b000110011;assign rom[7712] = 'b110000010;assign rom[7713] = 'b001101010;assign rom[7714] = 'b001011000;assign rom[7715] = 'b101001000;assign rom[7716] = 'b000101011;assign rom[7717] = 'b110000010;assign rom[7718] = 'b111000000;assign rom[7719] = 'b101001100;assign rom[7720] = 'b001001010;assign rom[7721] = 'b001000110;assign rom[7722] = 'b001100100;assign rom[7723] = 'b101100010;assign rom[7724] = 'b101001100;assign rom[7725] = 'b001001010;assign rom[7726] = 'b111011010;assign rom[7727] = 'b111011010;assign rom[7728] = 'b111011010;assign rom[7729] = 'b111011010;assign rom[7730] = 'b111011000;assign rom[7731] = 'b111011000;assign rom[7732] = 'b111011000;assign rom[7733] = 'b111011000;assign rom[7734] = 'b101111000;assign rom[7735] = 'b000110011;assign rom[7736] = 'b110000010;assign rom[7737] = 'b001101010;assign rom[7738] = 'b001011000;assign rom[7739] = 'b101001000;assign rom[7740] = 'b000101011;assign rom[7741] = 'b110000010;assign rom[7742] = 'b111000000;assign rom[7743] = 'b101001100;assign rom[7744] = 'b001001010;assign rom[7745] = 'b111111000;assign rom[7746] = 'b111101000;assign rom[7747] = 'b101001111;assign rom[7748] = 'b000111010;assign rom[7749] = 'b101110110;assign rom[7750] = 'b101100010;assign rom[7751] = 'b101001100;assign rom[7752] = 'b001001010;assign rom[7753] = 'b111011010;assign rom[7754] = 'b111011010;assign rom[7755] = 'b111011010;assign rom[7756] = 'b111011010;assign rom[7757] = 'b111011000;assign rom[7758] = 'b111011000;assign rom[7759] = 'b111011000;assign rom[7760] = 'b111011000;assign rom[7761] = 'b101111000;assign rom[7762] = 'b000110011;assign rom[7763] = 'b110000010;assign rom[7764] = 'b001101010;assign rom[7765] = 'b001011000;assign rom[7766] = 'b101001000;assign rom[7767] = 'b000101011;assign rom[7768] = 'b110000010;assign rom[7769] = 'b111000000;assign rom[7770] = 'b101001100;assign rom[7771] = 'b001001010;assign rom[7772] = 'b111111000;assign rom[7773] = 'b111101000;assign rom[7774] = 'b101001111;assign rom[7775] = 'b000111010;assign rom[7776] = 'b101110110;assign rom[7777] = 'b101100010;assign rom[7778] = 'b101001100;assign rom[7779] = 'b001001010;assign rom[7780] = 'b111011010;assign rom[7781] = 'b111011010;assign rom[7782] = 'b111011010;assign rom[7783] = 'b111011010;assign rom[7784] = 'b111011000;assign rom[7785] = 'b111011000;assign rom[7786] = 'b111011000;assign rom[7787] = 'b111011000;assign rom[7788] = 'b101111000;assign rom[7789] = 'b000110011;assign rom[7790] = 'b110000010;assign rom[7791] = 'b001101010;assign rom[7792] = 'b001011000;assign rom[7793] = 'b101001000;assign rom[7794] = 'b000101011;assign rom[7795] = 'b110000010;assign rom[7796] = 'b111000000;assign rom[7797] = 'b101001100;assign rom[7798] = 'b001001010;assign rom[7799] = 'b111111000;assign rom[7800] = 'b111101000;assign rom[7801] = 'b101001111;assign rom[7802] = 'b000111010;assign rom[7803] = 'b101110110;assign rom[7804] = 'b101100010;assign rom[7805] = 'b101001100;assign rom[7806] = 'b001001010;assign rom[7807] = 'b111011010;assign rom[7808] = 'b111011010;assign rom[7809] = 'b111011010;assign rom[7810] = 'b111011010;assign rom[7811] = 'b111011000;assign rom[7812] = 'b111011000;assign rom[7813] = 'b111011000;assign rom[7814] = 'b111011000;assign rom[7815] = 'b101111000;assign rom[7816] = 'b000110011;assign rom[7817] = 'b110000010;assign rom[7818] = 'b001101010;assign rom[7819] = 'b001011000;assign rom[7820] = 'b101001000;assign rom[7821] = 'b000101011;assign rom[7822] = 'b110000010;assign rom[7823] = 'b111000000;assign rom[7824] = 'b101001100;assign rom[7825] = 'b001001010;assign rom[7826] = 'b111111000;assign rom[7827] = 'b111101000;assign rom[7828] = 'b101001111;assign rom[7829] = 'b000111010;assign rom[7830] = 'b101110110;assign rom[7831] = 'b101100010;assign rom[7832] = 'b101001100;assign rom[7833] = 'b001001010;assign rom[7834] = 'b111011010;assign rom[7835] = 'b111011010;assign rom[7836] = 'b111011010;assign rom[7837] = 'b111011010;assign rom[7838] = 'b111011000;assign rom[7839] = 'b111011000;assign rom[7840] = 'b111011000;assign rom[7841] = 'b111011000;assign rom[7842] = 'b101111000;assign rom[7843] = 'b000110011;assign rom[7844] = 'b110000010;assign rom[7845] = 'b001101010;assign rom[7846] = 'b001011000;assign rom[7847] = 'b101001000;assign rom[7848] = 'b000101011;assign rom[7849] = 'b110000010;assign rom[7850] = 'b111000000;assign rom[7851] = 'b101001100;assign rom[7852] = 'b001001010;assign rom[7853] = 'b111111000;assign rom[7854] = 'b111101000;assign rom[7855] = 'b101001111;assign rom[7856] = 'b000111010;assign rom[7857] = 'b101110110;assign rom[7858] = 'b101100010;assign rom[7859] = 'b101001100;assign rom[7860] = 'b001001010;assign rom[7861] = 'b111011010;assign rom[7862] = 'b111011010;assign rom[7863] = 'b111011010;assign rom[7864] = 'b111011010;assign rom[7865] = 'b111011000;assign rom[7866] = 'b111011000;assign rom[7867] = 'b111011000;assign rom[7868] = 'b111011000;assign rom[7869] = 'b101111000;assign rom[7870] = 'b000110011;assign rom[7871] = 'b110000010;assign rom[7872] = 'b001101010;assign rom[7873] = 'b001011000;assign rom[7874] = 'b101001000;assign rom[7875] = 'b000101011;assign rom[7876] = 'b110000010;assign rom[7877] = 'b111000000;assign rom[7878] = 'b101001100;assign rom[7879] = 'b001001010;assign rom[7880] = 'b111111000;assign rom[7881] = 'b111101000;assign rom[7882] = 'b101001111;assign rom[7883] = 'b000111010;assign rom[7884] = 'b101110110;assign rom[7885] = 'b101100010;assign rom[7886] = 'b101001100;assign rom[7887] = 'b001001010;assign rom[7888] = 'b111011010;assign rom[7889] = 'b111011010;assign rom[7890] = 'b111011010;assign rom[7891] = 'b111011010;assign rom[7892] = 'b111011000;assign rom[7893] = 'b111011000;assign rom[7894] = 'b111011000;assign rom[7895] = 'b111011000;assign rom[7896] = 'b101111000;assign rom[7897] = 'b000110011;assign rom[7898] = 'b110000010;assign rom[7899] = 'b001101010;assign rom[7900] = 'b001011000;assign rom[7901] = 'b101001000;assign rom[7902] = 'b000101011;assign rom[7903] = 'b110000010;assign rom[7904] = 'b111000000;assign rom[7905] = 'b101001100;assign rom[7906] = 'b001001010;assign rom[7907] = 'b111111000;assign rom[7908] = 'b111101000;assign rom[7909] = 'b101001111;assign rom[7910] = 'b000111010;assign rom[7911] = 'b101110110;assign rom[7912] = 'b101100010;assign rom[7913] = 'b101001100;assign rom[7914] = 'b001001010;assign rom[7915] = 'b111011010;assign rom[7916] = 'b111011010;assign rom[7917] = 'b111011010;assign rom[7918] = 'b111011010;assign rom[7919] = 'b111011000;assign rom[7920] = 'b111011000;assign rom[7921] = 'b111011000;assign rom[7922] = 'b111011000;assign rom[7923] = 'b101111000;assign rom[7924] = 'b000110011;assign rom[7925] = 'b110000010;assign rom[7926] = 'b001101010;assign rom[7927] = 'b001011000;assign rom[7928] = 'b101001000;assign rom[7929] = 'b000101011;assign rom[7930] = 'b110000010;assign rom[7931] = 'b111000000;assign rom[7932] = 'b101001100;assign rom[7933] = 'b001001010;assign rom[7934] = 'b111111000;assign rom[7935] = 'b111101000;assign rom[7936] = 'b101001111;assign rom[7937] = 'b000111010;assign rom[7938] = 'b101110110;assign rom[7939] = 'b101100010;assign rom[7940] = 'b101001100;assign rom[7941] = 'b001001010;assign rom[7942] = 'b111011010;assign rom[7943] = 'b111011010;assign rom[7944] = 'b111011010;assign rom[7945] = 'b111011010;assign rom[7946] = 'b111011000;assign rom[7947] = 'b111011000;assign rom[7948] = 'b111011000;assign rom[7949] = 'b111011000;assign rom[7950] = 'b101111000;assign rom[7951] = 'b000110011;assign rom[7952] = 'b110000010;assign rom[7953] = 'b001101010;assign rom[7954] = 'b001011000;assign rom[7955] = 'b101001000;assign rom[7956] = 'b000101011;assign rom[7957] = 'b110000010;assign rom[7958] = 'b111000000;assign rom[7959] = 'b101001100;assign rom[7960] = 'b001001010;assign rom[7961] = 'b001000110;assign rom[7962] = 'b001100100;assign rom[7963] = 'b101100010;assign rom[7964] = 'b101001100;assign rom[7965] = 'b001001010;assign rom[7966] = 'b111011010;assign rom[7967] = 'b111011010;assign rom[7968] = 'b111011010;assign rom[7969] = 'b111011010;assign rom[7970] = 'b111011000;assign rom[7971] = 'b111011000;assign rom[7972] = 'b111011000;assign rom[7973] = 'b111011000;assign rom[7974] = 'b101111000;assign rom[7975] = 'b000110011;assign rom[7976] = 'b110000010;assign rom[7977] = 'b001101010;assign rom[7978] = 'b001011000;assign rom[7979] = 'b101001000;assign rom[7980] = 'b000101011;assign rom[7981] = 'b110000010;assign rom[7982] = 'b111000000;assign rom[7983] = 'b101001100;assign rom[7984] = 'b001001010;assign rom[7985] = 'b111111000;assign rom[7986] = 'b111101000;assign rom[7987] = 'b101001111;assign rom[7988] = 'b000111010;assign rom[7989] = 'b101110110;assign rom[7990] = 'b101100010;assign rom[7991] = 'b101001100;assign rom[7992] = 'b001001010;assign rom[7993] = 'b111011010;assign rom[7994] = 'b111011010;assign rom[7995] = 'b111011010;assign rom[7996] = 'b111011010;assign rom[7997] = 'b111011000;assign rom[7998] = 'b111011000;assign rom[7999] = 'b111011000;assign rom[8000] = 'b111011000;assign rom[8001] = 'b101111000;assign rom[8002] = 'b000110011;assign rom[8003] = 'b110000010;assign rom[8004] = 'b001101010;assign rom[8005] = 'b001011000;assign rom[8006] = 'b101001000;assign rom[8007] = 'b000101011;assign rom[8008] = 'b110000010;assign rom[8009] = 'b111000000;assign rom[8010] = 'b101001100;assign rom[8011] = 'b001001010;assign rom[8012] = 'b111111000;assign rom[8013] = 'b111101000;assign rom[8014] = 'b101001111;assign rom[8015] = 'b000111010;assign rom[8016] = 'b101110110;assign rom[8017] = 'b101100010;assign rom[8018] = 'b101001100;assign rom[8019] = 'b001001010;assign rom[8020] = 'b111011010;assign rom[8021] = 'b111011010;assign rom[8022] = 'b111011010;assign rom[8023] = 'b111011010;assign rom[8024] = 'b111011000;assign rom[8025] = 'b111011000;assign rom[8026] = 'b111011000;assign rom[8027] = 'b111011000;assign rom[8028] = 'b101111000;assign rom[8029] = 'b000110011;assign rom[8030] = 'b110000010;assign rom[8031] = 'b001101010;assign rom[8032] = 'b001011000;assign rom[8033] = 'b101001000;assign rom[8034] = 'b000101011;assign rom[8035] = 'b110000010;assign rom[8036] = 'b111000000;assign rom[8037] = 'b101001100;assign rom[8038] = 'b001001010;assign rom[8039] = 'b111111000;assign rom[8040] = 'b111101000;assign rom[8041] = 'b101001111;assign rom[8042] = 'b000111010;assign rom[8043] = 'b101110110;assign rom[8044] = 'b101100010;assign rom[8045] = 'b101001100;assign rom[8046] = 'b001001010;assign rom[8047] = 'b111011010;assign rom[8048] = 'b111011010;assign rom[8049] = 'b111011010;assign rom[8050] = 'b111011010;assign rom[8051] = 'b111011000;assign rom[8052] = 'b111011000;assign rom[8053] = 'b111011000;assign rom[8054] = 'b111011000;assign rom[8055] = 'b101111000;assign rom[8056] = 'b000110011;assign rom[8057] = 'b110000010;assign rom[8058] = 'b001101010;assign rom[8059] = 'b001011000;assign rom[8060] = 'b101001000;assign rom[8061] = 'b000101011;assign rom[8062] = 'b110000010;assign rom[8063] = 'b111000000;assign rom[8064] = 'b101001100;assign rom[8065] = 'b001001010;assign rom[8066] = 'b111111000;assign rom[8067] = 'b111101000;assign rom[8068] = 'b101001111;assign rom[8069] = 'b000111010;assign rom[8070] = 'b101110110;assign rom[8071] = 'b101100010;assign rom[8072] = 'b101001100;assign rom[8073] = 'b001001010;assign rom[8074] = 'b111011010;assign rom[8075] = 'b111011010;assign rom[8076] = 'b111011010;assign rom[8077] = 'b111011010;assign rom[8078] = 'b111011000;assign rom[8079] = 'b111011000;assign rom[8080] = 'b111011000;assign rom[8081] = 'b111011000;assign rom[8082] = 'b101111000;assign rom[8083] = 'b000110011;assign rom[8084] = 'b110000010;assign rom[8085] = 'b001101010;assign rom[8086] = 'b001011000;assign rom[8087] = 'b101001000;assign rom[8088] = 'b000101011;assign rom[8089] = 'b110000010;assign rom[8090] = 'b111000000;assign rom[8091] = 'b101001100;assign rom[8092] = 'b001001010;assign rom[8093] = 'b111111000;assign rom[8094] = 'b111101000;assign rom[8095] = 'b101001111;assign rom[8096] = 'b000111010;assign rom[8097] = 'b101110110;assign rom[8098] = 'b101100010;assign rom[8099] = 'b101001100;assign rom[8100] = 'b001001010;assign rom[8101] = 'b111011010;assign rom[8102] = 'b111011010;assign rom[8103] = 'b111011010;assign rom[8104] = 'b111011010;assign rom[8105] = 'b111011000;assign rom[8106] = 'b111011000;assign rom[8107] = 'b111011000;assign rom[8108] = 'b111011000;assign rom[8109] = 'b101111000;assign rom[8110] = 'b000110011;assign rom[8111] = 'b110000010;assign rom[8112] = 'b001101010;assign rom[8113] = 'b001011000;assign rom[8114] = 'b101001000;assign rom[8115] = 'b000101011;assign rom[8116] = 'b110000010;assign rom[8117] = 'b111000000;assign rom[8118] = 'b101001100;assign rom[8119] = 'b001001010;assign rom[8120] = 'b111111000;assign rom[8121] = 'b111101000;assign rom[8122] = 'b101001111;assign rom[8123] = 'b000111010;assign rom[8124] = 'b101110110;assign rom[8125] = 'b101100010;assign rom[8126] = 'b101001100;assign rom[8127] = 'b001001010;assign rom[8128] = 'b111011010;assign rom[8129] = 'b111011010;assign rom[8130] = 'b111011010;assign rom[8131] = 'b111011010;assign rom[8132] = 'b111011000;assign rom[8133] = 'b111011000;assign rom[8134] = 'b111011000;assign rom[8135] = 'b111011000;assign rom[8136] = 'b101111000;assign rom[8137] = 'b000110011;assign rom[8138] = 'b110000010;assign rom[8139] = 'b001101010;assign rom[8140] = 'b001011000;assign rom[8141] = 'b101001000;assign rom[8142] = 'b000101011;assign rom[8143] = 'b110000010;assign rom[8144] = 'b111000000;assign rom[8145] = 'b101001100;assign rom[8146] = 'b001001010;assign rom[8147] = 'b111111000;assign rom[8148] = 'b111101000;assign rom[8149] = 'b101001111;assign rom[8150] = 'b000111010;assign rom[8151] = 'b101110110;assign rom[8152] = 'b101100010;assign rom[8153] = 'b101001100;assign rom[8154] = 'b001001010;assign rom[8155] = 'b111011010;assign rom[8156] = 'b111011010;assign rom[8157] = 'b111011010;assign rom[8158] = 'b111011010;assign rom[8159] = 'b111011000;assign rom[8160] = 'b111011000;assign rom[8161] = 'b111011000;assign rom[8162] = 'b111011000;assign rom[8163] = 'b101111000;assign rom[8164] = 'b000110011;assign rom[8165] = 'b110000010;assign rom[8166] = 'b001101010;assign rom[8167] = 'b001011000;assign rom[8168] = 'b101001000;assign rom[8169] = 'b000101011;assign rom[8170] = 'b110000010;assign rom[8171] = 'b111000000;assign rom[8172] = 'b101001100;assign rom[8173] = 'b001001010;assign rom[8174] = 'b111111000;assign rom[8175] = 'b111101000;assign rom[8176] = 'b101001111;assign rom[8177] = 'b000111010;assign rom[8178] = 'b101110110;assign rom[8179] = 'b101100010;assign rom[8180] = 'b101001100;assign rom[8181] = 'b001001010;assign rom[8182] = 'b111011010;assign rom[8183] = 'b111011010;assign rom[8184] = 'b111011010;assign rom[8185] = 'b111011010;assign rom[8186] = 'b111011000;assign rom[8187] = 'b111011000;assign rom[8188] = 'b111011000;assign rom[8189] = 'b111011000;assign rom[8190] = 'b101111000;assign rom[8191] = 'b000110011;assign rom[8192] = 'b110000010;assign rom[8193] = 'b001101010;assign rom[8194] = 'b001011000;assign rom[8195] = 'b101001000;assign rom[8196] = 'b000101011;assign rom[8197] = 'b110000010;assign rom[8198] = 'b111000000;assign rom[8199] = 'b101001100;assign rom[8200] = 'b001001010;assign rom[8201] = 'b001000110;assign rom[8202] = 'b001100100;assign rom[8203] = 'b101100010;assign rom[8204] = 'b101001100;assign rom[8205] = 'b001001010;assign rom[8206] = 'b111011010;assign rom[8207] = 'b111011010;assign rom[8208] = 'b111011010;assign rom[8209] = 'b111011010;assign rom[8210] = 'b111011000;assign rom[8211] = 'b111011000;assign rom[8212] = 'b111011000;assign rom[8213] = 'b111011000;assign rom[8214] = 'b101111000;assign rom[8215] = 'b000110011;assign rom[8216] = 'b110000010;assign rom[8217] = 'b001101010;assign rom[8218] = 'b001011000;assign rom[8219] = 'b101001000;assign rom[8220] = 'b000101011;assign rom[8221] = 'b110000010;assign rom[8222] = 'b111000000;assign rom[8223] = 'b101001100;assign rom[8224] = 'b001001010;assign rom[8225] = 'b111111000;assign rom[8226] = 'b111101000;assign rom[8227] = 'b101001111;assign rom[8228] = 'b000111010;assign rom[8229] = 'b101110110;assign rom[8230] = 'b101100010;assign rom[8231] = 'b101001100;assign rom[8232] = 'b001001010;assign rom[8233] = 'b111011010;assign rom[8234] = 'b111011010;assign rom[8235] = 'b111011010;assign rom[8236] = 'b111011010;assign rom[8237] = 'b111011000;assign rom[8238] = 'b111011000;assign rom[8239] = 'b111011000;assign rom[8240] = 'b111011000;assign rom[8241] = 'b101111000;assign rom[8242] = 'b000110011;assign rom[8243] = 'b110000010;assign rom[8244] = 'b001101010;assign rom[8245] = 'b001011000;assign rom[8246] = 'b101001000;assign rom[8247] = 'b000101011;assign rom[8248] = 'b110000010;assign rom[8249] = 'b111000000;assign rom[8250] = 'b101001100;assign rom[8251] = 'b001001010;assign rom[8252] = 'b111111000;assign rom[8253] = 'b111101000;assign rom[8254] = 'b101001111;assign rom[8255] = 'b000111010;assign rom[8256] = 'b101110110;assign rom[8257] = 'b101100010;assign rom[8258] = 'b101001100;assign rom[8259] = 'b001001010;assign rom[8260] = 'b111011010;assign rom[8261] = 'b111011010;assign rom[8262] = 'b111011010;assign rom[8263] = 'b111011010;assign rom[8264] = 'b111011000;assign rom[8265] = 'b111011000;assign rom[8266] = 'b111011000;assign rom[8267] = 'b111011000;assign rom[8268] = 'b101111000;assign rom[8269] = 'b000110011;assign rom[8270] = 'b110000010;assign rom[8271] = 'b001101010;assign rom[8272] = 'b001011000;assign rom[8273] = 'b101001000;assign rom[8274] = 'b000101011;assign rom[8275] = 'b110000010;assign rom[8276] = 'b111000000;assign rom[8277] = 'b101001100;assign rom[8278] = 'b001001010;assign rom[8279] = 'b111111000;assign rom[8280] = 'b111101000;assign rom[8281] = 'b101001111;assign rom[8282] = 'b000111010;assign rom[8283] = 'b101110110;assign rom[8284] = 'b101100010;assign rom[8285] = 'b101001100;assign rom[8286] = 'b001001010;assign rom[8287] = 'b111011010;assign rom[8288] = 'b111011010;assign rom[8289] = 'b111011010;assign rom[8290] = 'b111011010;assign rom[8291] = 'b111011000;assign rom[8292] = 'b111011000;assign rom[8293] = 'b111011000;assign rom[8294] = 'b111011000;assign rom[8295] = 'b101111000;assign rom[8296] = 'b000110011;assign rom[8297] = 'b110000010;assign rom[8298] = 'b001101010;assign rom[8299] = 'b001011000;assign rom[8300] = 'b101001000;assign rom[8301] = 'b000101011;assign rom[8302] = 'b110000010;assign rom[8303] = 'b111000000;assign rom[8304] = 'b101001100;assign rom[8305] = 'b001001010;assign rom[8306] = 'b111111000;assign rom[8307] = 'b111101000;assign rom[8308] = 'b101001111;assign rom[8309] = 'b000111010;assign rom[8310] = 'b101110110;assign rom[8311] = 'b101100010;assign rom[8312] = 'b101001100;assign rom[8313] = 'b001001010;assign rom[8314] = 'b111011010;assign rom[8315] = 'b111011010;assign rom[8316] = 'b111011010;assign rom[8317] = 'b111011010;assign rom[8318] = 'b111011000;assign rom[8319] = 'b111011000;assign rom[8320] = 'b111011000;assign rom[8321] = 'b111011000;assign rom[8322] = 'b101111000;assign rom[8323] = 'b000110011;assign rom[8324] = 'b110000010;assign rom[8325] = 'b001101010;assign rom[8326] = 'b001011000;assign rom[8327] = 'b101001000;assign rom[8328] = 'b000101011;assign rom[8329] = 'b110000010;assign rom[8330] = 'b111000000;assign rom[8331] = 'b101001100;assign rom[8332] = 'b001001010;assign rom[8333] = 'b111111000;assign rom[8334] = 'b111101000;assign rom[8335] = 'b101001111;assign rom[8336] = 'b000111010;assign rom[8337] = 'b101110110;assign rom[8338] = 'b101100010;assign rom[8339] = 'b101001100;assign rom[8340] = 'b001001010;assign rom[8341] = 'b111011010;assign rom[8342] = 'b111011010;assign rom[8343] = 'b111011010;assign rom[8344] = 'b111011010;assign rom[8345] = 'b111011000;assign rom[8346] = 'b111011000;assign rom[8347] = 'b111011000;assign rom[8348] = 'b111011000;assign rom[8349] = 'b101111000;assign rom[8350] = 'b000110011;assign rom[8351] = 'b110000010;assign rom[8352] = 'b001101010;assign rom[8353] = 'b001011000;assign rom[8354] = 'b101001000;assign rom[8355] = 'b000101011;assign rom[8356] = 'b110000010;assign rom[8357] = 'b111000000;assign rom[8358] = 'b101001100;assign rom[8359] = 'b001001010;assign rom[8360] = 'b111111000;assign rom[8361] = 'b111101000;assign rom[8362] = 'b101001111;assign rom[8363] = 'b000111010;assign rom[8364] = 'b101110110;assign rom[8365] = 'b101100010;assign rom[8366] = 'b101001100;assign rom[8367] = 'b001001010;assign rom[8368] = 'b111011010;assign rom[8369] = 'b111011010;assign rom[8370] = 'b111011010;assign rom[8371] = 'b111011010;assign rom[8372] = 'b111011000;assign rom[8373] = 'b111011000;assign rom[8374] = 'b111011000;assign rom[8375] = 'b111011000;assign rom[8376] = 'b101111000;assign rom[8377] = 'b000110011;assign rom[8378] = 'b110000010;assign rom[8379] = 'b001101010;assign rom[8380] = 'b001011000;assign rom[8381] = 'b101001000;assign rom[8382] = 'b000101011;assign rom[8383] = 'b110000010;assign rom[8384] = 'b111000000;assign rom[8385] = 'b101001100;assign rom[8386] = 'b001001010;assign rom[8387] = 'b111111000;assign rom[8388] = 'b111101000;assign rom[8389] = 'b101001111;assign rom[8390] = 'b000111010;assign rom[8391] = 'b101110110;assign rom[8392] = 'b101100010;assign rom[8393] = 'b101001100;assign rom[8394] = 'b001001010;assign rom[8395] = 'b111011010;assign rom[8396] = 'b111011010;assign rom[8397] = 'b111011010;assign rom[8398] = 'b111011010;assign rom[8399] = 'b111011000;assign rom[8400] = 'b111011000;assign rom[8401] = 'b111011000;assign rom[8402] = 'b111011000;assign rom[8403] = 'b101111000;assign rom[8404] = 'b000110011;assign rom[8405] = 'b110000010;assign rom[8406] = 'b001101010;assign rom[8407] = 'b001011000;assign rom[8408] = 'b101001000;assign rom[8409] = 'b000101011;assign rom[8410] = 'b110000010;assign rom[8411] = 'b111000000;assign rom[8412] = 'b101001100;assign rom[8413] = 'b001001010;assign rom[8414] = 'b111111000;assign rom[8415] = 'b111101000;assign rom[8416] = 'b101001111;assign rom[8417] = 'b000111010;assign rom[8418] = 'b101110110;assign rom[8419] = 'b101100010;assign rom[8420] = 'b101001100;assign rom[8421] = 'b001001010;assign rom[8422] = 'b111011010;assign rom[8423] = 'b111011010;assign rom[8424] = 'b111011010;assign rom[8425] = 'b111011010;assign rom[8426] = 'b111011000;assign rom[8427] = 'b111011000;assign rom[8428] = 'b111011000;assign rom[8429] = 'b111011000;assign rom[8430] = 'b101111000;assign rom[8431] = 'b000110011;assign rom[8432] = 'b110000010;assign rom[8433] = 'b001101010;assign rom[8434] = 'b001011000;assign rom[8435] = 'b101001000;assign rom[8436] = 'b000101011;assign rom[8437] = 'b110000010;assign rom[8438] = 'b111000000;assign rom[8439] = 'b101001100;assign rom[8440] = 'b001001010;assign rom[8441] = 'b001000110;assign rom[8442] = 'b001100100;assign rom[8443] = 'b101100010;assign rom[8444] = 'b101001100;assign rom[8445] = 'b001001010;assign rom[8446] = 'b111011010;assign rom[8447] = 'b111011010;assign rom[8448] = 'b111011010;assign rom[8449] = 'b111011010;assign rom[8450] = 'b111011000;assign rom[8451] = 'b111011000;assign rom[8452] = 'b111011000;assign rom[8453] = 'b111011000;assign rom[8454] = 'b101111000;assign rom[8455] = 'b000110011;assign rom[8456] = 'b110000010;assign rom[8457] = 'b001101010;assign rom[8458] = 'b001011000;assign rom[8459] = 'b101001000;assign rom[8460] = 'b000101011;assign rom[8461] = 'b110000010;assign rom[8462] = 'b111000000;assign rom[8463] = 'b101001100;assign rom[8464] = 'b001001010;assign rom[8465] = 'b111111000;assign rom[8466] = 'b111101000;assign rom[8467] = 'b101001111;assign rom[8468] = 'b000111010;assign rom[8469] = 'b101110110;assign rom[8470] = 'b101100010;assign rom[8471] = 'b101001100;assign rom[8472] = 'b001001010;assign rom[8473] = 'b111011010;assign rom[8474] = 'b111011010;assign rom[8475] = 'b111011010;assign rom[8476] = 'b111011010;assign rom[8477] = 'b111011000;assign rom[8478] = 'b111011000;assign rom[8479] = 'b111011000;assign rom[8480] = 'b111011000;assign rom[8481] = 'b101111000;assign rom[8482] = 'b000110011;assign rom[8483] = 'b110000010;assign rom[8484] = 'b001101010;assign rom[8485] = 'b001011000;assign rom[8486] = 'b101001000;assign rom[8487] = 'b000101011;assign rom[8488] = 'b110000010;assign rom[8489] = 'b111000000;assign rom[8490] = 'b101001100;assign rom[8491] = 'b001001010;assign rom[8492] = 'b111111000;assign rom[8493] = 'b111101000;assign rom[8494] = 'b101001111;assign rom[8495] = 'b000111010;assign rom[8496] = 'b101110110;assign rom[8497] = 'b101100010;assign rom[8498] = 'b101001100;assign rom[8499] = 'b001001010;assign rom[8500] = 'b111011010;assign rom[8501] = 'b111011010;assign rom[8502] = 'b111011010;assign rom[8503] = 'b111011010;assign rom[8504] = 'b111011000;assign rom[8505] = 'b111011000;assign rom[8506] = 'b111011000;assign rom[8507] = 'b111011000;assign rom[8508] = 'b101111000;assign rom[8509] = 'b000110011;assign rom[8510] = 'b110000010;assign rom[8511] = 'b001101010;assign rom[8512] = 'b001011000;assign rom[8513] = 'b101001000;assign rom[8514] = 'b000101011;assign rom[8515] = 'b110000010;assign rom[8516] = 'b111000000;assign rom[8517] = 'b101001100;assign rom[8518] = 'b001001010;assign rom[8519] = 'b111111000;assign rom[8520] = 'b111101000;assign rom[8521] = 'b101001111;assign rom[8522] = 'b000111010;assign rom[8523] = 'b101110110;assign rom[8524] = 'b101100010;assign rom[8525] = 'b101001100;assign rom[8526] = 'b001001010;assign rom[8527] = 'b111011010;assign rom[8528] = 'b111011010;assign rom[8529] = 'b111011010;assign rom[8530] = 'b111011010;assign rom[8531] = 'b111011000;assign rom[8532] = 'b111011000;assign rom[8533] = 'b111011000;assign rom[8534] = 'b111011000;assign rom[8535] = 'b101111000;assign rom[8536] = 'b000110011;assign rom[8537] = 'b110000010;assign rom[8538] = 'b001101010;assign rom[8539] = 'b001011000;assign rom[8540] = 'b101001000;assign rom[8541] = 'b000101011;assign rom[8542] = 'b110000010;assign rom[8543] = 'b111000000;assign rom[8544] = 'b101001100;assign rom[8545] = 'b001001010;assign rom[8546] = 'b111111000;assign rom[8547] = 'b111101000;assign rom[8548] = 'b101001111;assign rom[8549] = 'b000111010;assign rom[8550] = 'b101110110;assign rom[8551] = 'b101100010;assign rom[8552] = 'b101001100;assign rom[8553] = 'b001001010;assign rom[8554] = 'b111011010;assign rom[8555] = 'b111011010;assign rom[8556] = 'b111011010;assign rom[8557] = 'b111011010;assign rom[8558] = 'b111011000;assign rom[8559] = 'b111011000;assign rom[8560] = 'b111011000;assign rom[8561] = 'b111011000;assign rom[8562] = 'b101111000;assign rom[8563] = 'b000110011;assign rom[8564] = 'b110000010;assign rom[8565] = 'b001101010;assign rom[8566] = 'b001011000;assign rom[8567] = 'b101001000;assign rom[8568] = 'b000101011;assign rom[8569] = 'b110000010;assign rom[8570] = 'b111000000;assign rom[8571] = 'b101001100;assign rom[8572] = 'b001001010;assign rom[8573] = 'b111111000;assign rom[8574] = 'b111101000;assign rom[8575] = 'b101001111;assign rom[8576] = 'b000111010;assign rom[8577] = 'b101110110;assign rom[8578] = 'b101100010;assign rom[8579] = 'b101001100;assign rom[8580] = 'b001001010;assign rom[8581] = 'b111011010;assign rom[8582] = 'b111011010;assign rom[8583] = 'b111011010;assign rom[8584] = 'b111011010;assign rom[8585] = 'b111011000;assign rom[8586] = 'b111011000;assign rom[8587] = 'b111011000;assign rom[8588] = 'b111011000;assign rom[8589] = 'b101111000;assign rom[8590] = 'b000110011;assign rom[8591] = 'b110000010;assign rom[8592] = 'b001101010;assign rom[8593] = 'b001011000;assign rom[8594] = 'b101001000;assign rom[8595] = 'b000101011;assign rom[8596] = 'b110000010;assign rom[8597] = 'b111000000;assign rom[8598] = 'b101001100;assign rom[8599] = 'b001001010;assign rom[8600] = 'b111111000;assign rom[8601] = 'b111101000;assign rom[8602] = 'b101001111;assign rom[8603] = 'b000111010;assign rom[8604] = 'b101110110;assign rom[8605] = 'b101100010;assign rom[8606] = 'b101001100;assign rom[8607] = 'b001001010;assign rom[8608] = 'b111011010;assign rom[8609] = 'b111011010;assign rom[8610] = 'b111011010;assign rom[8611] = 'b111011010;assign rom[8612] = 'b111011000;assign rom[8613] = 'b111011000;assign rom[8614] = 'b111011000;assign rom[8615] = 'b111011000;assign rom[8616] = 'b101111000;assign rom[8617] = 'b000110011;assign rom[8618] = 'b110000010;assign rom[8619] = 'b001101010;assign rom[8620] = 'b001011000;assign rom[8621] = 'b101001000;assign rom[8622] = 'b000101011;assign rom[8623] = 'b110000010;assign rom[8624] = 'b111000000;assign rom[8625] = 'b101001100;assign rom[8626] = 'b001001010;assign rom[8627] = 'b111111000;assign rom[8628] = 'b111101000;assign rom[8629] = 'b101001111;assign rom[8630] = 'b000111010;assign rom[8631] = 'b101110110;assign rom[8632] = 'b101100010;assign rom[8633] = 'b101001100;assign rom[8634] = 'b001001010;assign rom[8635] = 'b111011010;assign rom[8636] = 'b111011010;assign rom[8637] = 'b111011010;assign rom[8638] = 'b111011010;assign rom[8639] = 'b111011000;assign rom[8640] = 'b111011000;assign rom[8641] = 'b111011000;assign rom[8642] = 'b111011000;assign rom[8643] = 'b101111000;assign rom[8644] = 'b000110011;assign rom[8645] = 'b110000010;assign rom[8646] = 'b001101010;assign rom[8647] = 'b001011000;assign rom[8648] = 'b101001000;assign rom[8649] = 'b000101011;assign rom[8650] = 'b110000010;assign rom[8651] = 'b111000000;assign rom[8652] = 'b101001100;assign rom[8653] = 'b001001010;assign rom[8654] = 'b111111000;assign rom[8655] = 'b111101000;assign rom[8656] = 'b101001111;assign rom[8657] = 'b000111010;assign rom[8658] = 'b101110110;assign rom[8659] = 'b101100010;assign rom[8660] = 'b101001100;assign rom[8661] = 'b001001010;assign rom[8662] = 'b111011010;assign rom[8663] = 'b111011010;assign rom[8664] = 'b111011010;assign rom[8665] = 'b111011010;assign rom[8666] = 'b111011000;assign rom[8667] = 'b111011000;assign rom[8668] = 'b111011000;assign rom[8669] = 'b111011000;assign rom[8670] = 'b101111000;assign rom[8671] = 'b000110011;assign rom[8672] = 'b110000010;assign rom[8673] = 'b001101010;assign rom[8674] = 'b001011000;assign rom[8675] = 'b101001000;assign rom[8676] = 'b000101011;assign rom[8677] = 'b110000010;assign rom[8678] = 'b111000000;assign rom[8679] = 'b101001100;assign rom[8680] = 'b001001010;assign rom[8681] = 'b001000110;assign rom[8682] = 'b001100100;assign rom[8683] = 'b101100010;assign rom[8684] = 'b101001100;assign rom[8685] = 'b001001010;assign rom[8686] = 'b111011010;assign rom[8687] = 'b111011010;assign rom[8688] = 'b111011010;assign rom[8689] = 'b111011010;assign rom[8690] = 'b111011000;assign rom[8691] = 'b111011000;assign rom[8692] = 'b111011000;assign rom[8693] = 'b111011000;assign rom[8694] = 'b101111000;assign rom[8695] = 'b000110011;assign rom[8696] = 'b110000010;assign rom[8697] = 'b001101010;assign rom[8698] = 'b001011000;assign rom[8699] = 'b101001000;assign rom[8700] = 'b000101011;assign rom[8701] = 'b110000010;assign rom[8702] = 'b111000000;assign rom[8703] = 'b101001100;assign rom[8704] = 'b001001010;assign rom[8705] = 'b111111000;assign rom[8706] = 'b111101000;assign rom[8707] = 'b101001111;assign rom[8708] = 'b000111010;assign rom[8709] = 'b101110110;assign rom[8710] = 'b101100010;assign rom[8711] = 'b101001100;assign rom[8712] = 'b001001010;assign rom[8713] = 'b111011010;assign rom[8714] = 'b111011010;assign rom[8715] = 'b111011010;assign rom[8716] = 'b111011010;assign rom[8717] = 'b111011000;assign rom[8718] = 'b111011000;assign rom[8719] = 'b111011000;assign rom[8720] = 'b111011000;assign rom[8721] = 'b101111000;assign rom[8722] = 'b000110011;assign rom[8723] = 'b110000010;assign rom[8724] = 'b001101010;assign rom[8725] = 'b001011000;assign rom[8726] = 'b101001000;assign rom[8727] = 'b000101011;assign rom[8728] = 'b110000010;assign rom[8729] = 'b111000000;assign rom[8730] = 'b101001100;assign rom[8731] = 'b001001010;assign rom[8732] = 'b111111000;assign rom[8733] = 'b111101000;assign rom[8734] = 'b101001111;assign rom[8735] = 'b000111010;assign rom[8736] = 'b101110110;assign rom[8737] = 'b101100010;assign rom[8738] = 'b101001100;assign rom[8739] = 'b001001010;assign rom[8740] = 'b111011010;assign rom[8741] = 'b111011010;assign rom[8742] = 'b111011010;assign rom[8743] = 'b111011010;assign rom[8744] = 'b111011000;assign rom[8745] = 'b111011000;assign rom[8746] = 'b111011000;assign rom[8747] = 'b111011000;assign rom[8748] = 'b101111000;assign rom[8749] = 'b000110011;assign rom[8750] = 'b110000010;assign rom[8751] = 'b001101010;assign rom[8752] = 'b001011000;assign rom[8753] = 'b101001000;assign rom[8754] = 'b000101011;assign rom[8755] = 'b110000010;assign rom[8756] = 'b111000000;assign rom[8757] = 'b101001100;assign rom[8758] = 'b001001010;assign rom[8759] = 'b111111000;assign rom[8760] = 'b111101000;assign rom[8761] = 'b101001111;assign rom[8762] = 'b000111010;assign rom[8763] = 'b101110110;assign rom[8764] = 'b101100010;assign rom[8765] = 'b101001100;assign rom[8766] = 'b001001010;assign rom[8767] = 'b111011010;assign rom[8768] = 'b111011010;assign rom[8769] = 'b111011010;assign rom[8770] = 'b111011010;assign rom[8771] = 'b111011000;assign rom[8772] = 'b111011000;assign rom[8773] = 'b111011000;assign rom[8774] = 'b111011000;assign rom[8775] = 'b101111000;assign rom[8776] = 'b000110011;assign rom[8777] = 'b110000010;assign rom[8778] = 'b001101010;assign rom[8779] = 'b001011000;assign rom[8780] = 'b101001000;assign rom[8781] = 'b000101011;assign rom[8782] = 'b110000010;assign rom[8783] = 'b111000000;assign rom[8784] = 'b101001100;assign rom[8785] = 'b001001010;assign rom[8786] = 'b111111000;assign rom[8787] = 'b111101000;assign rom[8788] = 'b101001111;assign rom[8789] = 'b000111010;assign rom[8790] = 'b101110110;assign rom[8791] = 'b101100010;assign rom[8792] = 'b101001100;assign rom[8793] = 'b001001010;assign rom[8794] = 'b111011010;assign rom[8795] = 'b111011010;assign rom[8796] = 'b111011010;assign rom[8797] = 'b111011010;assign rom[8798] = 'b111011000;assign rom[8799] = 'b111011000;assign rom[8800] = 'b111011000;assign rom[8801] = 'b111011000;assign rom[8802] = 'b101111000;assign rom[8803] = 'b000110011;assign rom[8804] = 'b110000010;assign rom[8805] = 'b001101010;assign rom[8806] = 'b001011000;assign rom[8807] = 'b101001000;assign rom[8808] = 'b000101011;assign rom[8809] = 'b110000010;assign rom[8810] = 'b111000000;assign rom[8811] = 'b101001100;assign rom[8812] = 'b001001010;assign rom[8813] = 'b111111000;assign rom[8814] = 'b111101000;assign rom[8815] = 'b101001111;assign rom[8816] = 'b000111010;assign rom[8817] = 'b101110110;assign rom[8818] = 'b101100010;assign rom[8819] = 'b101001100;assign rom[8820] = 'b001001010;assign rom[8821] = 'b111011010;assign rom[8822] = 'b111011010;assign rom[8823] = 'b111011010;assign rom[8824] = 'b111011010;assign rom[8825] = 'b111011000;assign rom[8826] = 'b111011000;assign rom[8827] = 'b111011000;assign rom[8828] = 'b111011000;assign rom[8829] = 'b101111000;assign rom[8830] = 'b000110011;assign rom[8831] = 'b110000010;assign rom[8832] = 'b001101010;assign rom[8833] = 'b001011000;assign rom[8834] = 'b101001000;assign rom[8835] = 'b000101011;assign rom[8836] = 'b110000010;assign rom[8837] = 'b111000000;assign rom[8838] = 'b101001100;assign rom[8839] = 'b001001010;assign rom[8840] = 'b111111000;assign rom[8841] = 'b111101000;assign rom[8842] = 'b101001111;assign rom[8843] = 'b000111010;assign rom[8844] = 'b101110110;assign rom[8845] = 'b101100010;assign rom[8846] = 'b101001100;assign rom[8847] = 'b001001010;assign rom[8848] = 'b111011010;assign rom[8849] = 'b111011010;assign rom[8850] = 'b111011010;assign rom[8851] = 'b111011010;assign rom[8852] = 'b111011000;assign rom[8853] = 'b111011000;assign rom[8854] = 'b111011000;assign rom[8855] = 'b111011000;assign rom[8856] = 'b101111000;assign rom[8857] = 'b000110011;assign rom[8858] = 'b110000010;assign rom[8859] = 'b001101010;assign rom[8860] = 'b001011000;assign rom[8861] = 'b101001000;assign rom[8862] = 'b000101011;assign rom[8863] = 'b110000010;assign rom[8864] = 'b111000000;assign rom[8865] = 'b101001100;assign rom[8866] = 'b001001010;assign rom[8867] = 'b111111000;assign rom[8868] = 'b111101000;assign rom[8869] = 'b101001111;assign rom[8870] = 'b000111010;assign rom[8871] = 'b101110110;assign rom[8872] = 'b101100010;assign rom[8873] = 'b101001100;assign rom[8874] = 'b001001010;assign rom[8875] = 'b111011010;assign rom[8876] = 'b111011010;assign rom[8877] = 'b111011010;assign rom[8878] = 'b111011010;assign rom[8879] = 'b111011000;assign rom[8880] = 'b111011000;assign rom[8881] = 'b111011000;assign rom[8882] = 'b111011000;assign rom[8883] = 'b101111000;assign rom[8884] = 'b000110011;assign rom[8885] = 'b110000010;assign rom[8886] = 'b001101010;assign rom[8887] = 'b001011000;assign rom[8888] = 'b101001000;assign rom[8889] = 'b000101011;assign rom[8890] = 'b110000010;assign rom[8891] = 'b111000000;assign rom[8892] = 'b101001100;assign rom[8893] = 'b001001010;assign rom[8894] = 'b111111000;assign rom[8895] = 'b111101000;assign rom[8896] = 'b101001111;assign rom[8897] = 'b000111010;assign rom[8898] = 'b101110110;assign rom[8899] = 'b101100010;assign rom[8900] = 'b101001100;assign rom[8901] = 'b001001010;assign rom[8902] = 'b111011010;assign rom[8903] = 'b111011010;assign rom[8904] = 'b111011010;assign rom[8905] = 'b111011010;assign rom[8906] = 'b111011000;assign rom[8907] = 'b111011000;assign rom[8908] = 'b111011000;assign rom[8909] = 'b111011000;assign rom[8910] = 'b101111000;assign rom[8911] = 'b000110011;assign rom[8912] = 'b110000010;assign rom[8913] = 'b001101010;assign rom[8914] = 'b001011000;assign rom[8915] = 'b101001000;assign rom[8916] = 'b000101011;assign rom[8917] = 'b110000010;assign rom[8918] = 'b111000000;assign rom[8919] = 'b101001100;assign rom[8920] = 'b001001010;assign rom[8921] = 'b001000110;assign rom[8922] = 'b001100100;assign rom[8923] = 'b101100010;assign rom[8924] = 'b101001100;assign rom[8925] = 'b001001010;assign rom[8926] = 'b111011010;assign rom[8927] = 'b111011010;assign rom[8928] = 'b111011010;assign rom[8929] = 'b111011010;assign rom[8930] = 'b111011000;assign rom[8931] = 'b111011000;assign rom[8932] = 'b111011000;assign rom[8933] = 'b111011000;assign rom[8934] = 'b101111000;assign rom[8935] = 'b000110011;assign rom[8936] = 'b110000010;assign rom[8937] = 'b001101010;assign rom[8938] = 'b001011000;assign rom[8939] = 'b101001000;assign rom[8940] = 'b000101011;assign rom[8941] = 'b110000010;assign rom[8942] = 'b111000000;assign rom[8943] = 'b101001100;assign rom[8944] = 'b001001010;assign rom[8945] = 'b111111000;assign rom[8946] = 'b111101000;assign rom[8947] = 'b101001111;assign rom[8948] = 'b000111010;assign rom[8949] = 'b101110110;assign rom[8950] = 'b101100010;assign rom[8951] = 'b101001100;assign rom[8952] = 'b001001010;assign rom[8953] = 'b111011010;assign rom[8954] = 'b111011010;assign rom[8955] = 'b111011010;assign rom[8956] = 'b111011010;assign rom[8957] = 'b111011000;assign rom[8958] = 'b111011000;assign rom[8959] = 'b111011000;assign rom[8960] = 'b111011000;assign rom[8961] = 'b101111000;assign rom[8962] = 'b000110011;assign rom[8963] = 'b110000010;assign rom[8964] = 'b001101010;assign rom[8965] = 'b001011000;assign rom[8966] = 'b101001000;assign rom[8967] = 'b000101011;assign rom[8968] = 'b110000010;assign rom[8969] = 'b111000000;assign rom[8970] = 'b101001100;assign rom[8971] = 'b001001010;assign rom[8972] = 'b111111000;assign rom[8973] = 'b111101000;assign rom[8974] = 'b101001111;assign rom[8975] = 'b000111010;assign rom[8976] = 'b101110110;assign rom[8977] = 'b101100010;assign rom[8978] = 'b101001100;assign rom[8979] = 'b001001010;assign rom[8980] = 'b111011010;assign rom[8981] = 'b111011010;assign rom[8982] = 'b111011010;assign rom[8983] = 'b111011010;assign rom[8984] = 'b111011000;assign rom[8985] = 'b111011000;assign rom[8986] = 'b111011000;assign rom[8987] = 'b111011000;assign rom[8988] = 'b101111000;assign rom[8989] = 'b000110011;assign rom[8990] = 'b110000010;assign rom[8991] = 'b001101010;assign rom[8992] = 'b001011000;assign rom[8993] = 'b101001000;assign rom[8994] = 'b000101011;assign rom[8995] = 'b110000010;assign rom[8996] = 'b111000000;assign rom[8997] = 'b101001100;assign rom[8998] = 'b001001010;assign rom[8999] = 'b111111000;assign rom[9000] = 'b111101000;assign rom[9001] = 'b101001111;assign rom[9002] = 'b000111010;assign rom[9003] = 'b101110110;assign rom[9004] = 'b101100010;assign rom[9005] = 'b101001100;assign rom[9006] = 'b001001010;assign rom[9007] = 'b111011010;assign rom[9008] = 'b111011010;assign rom[9009] = 'b111011010;assign rom[9010] = 'b111011010;assign rom[9011] = 'b111011000;assign rom[9012] = 'b111011000;assign rom[9013] = 'b111011000;assign rom[9014] = 'b111011000;assign rom[9015] = 'b101111000;assign rom[9016] = 'b000110011;assign rom[9017] = 'b110000010;assign rom[9018] = 'b001101010;assign rom[9019] = 'b001011000;assign rom[9020] = 'b101001000;assign rom[9021] = 'b000101011;assign rom[9022] = 'b110000010;assign rom[9023] = 'b111000000;assign rom[9024] = 'b101001100;assign rom[9025] = 'b001001010;assign rom[9026] = 'b111111000;assign rom[9027] = 'b111101000;assign rom[9028] = 'b101001111;assign rom[9029] = 'b000111010;assign rom[9030] = 'b101110110;assign rom[9031] = 'b101100010;assign rom[9032] = 'b101001100;assign rom[9033] = 'b001001010;assign rom[9034] = 'b111011010;assign rom[9035] = 'b111011010;assign rom[9036] = 'b111011010;assign rom[9037] = 'b111011010;assign rom[9038] = 'b111011000;assign rom[9039] = 'b111011000;assign rom[9040] = 'b111011000;assign rom[9041] = 'b111011000;assign rom[9042] = 'b101111000;assign rom[9043] = 'b000110011;assign rom[9044] = 'b110000010;assign rom[9045] = 'b001101010;assign rom[9046] = 'b001011000;assign rom[9047] = 'b101001000;assign rom[9048] = 'b000101011;assign rom[9049] = 'b110000010;assign rom[9050] = 'b111000000;assign rom[9051] = 'b101001100;assign rom[9052] = 'b001001010;assign rom[9053] = 'b111111000;assign rom[9054] = 'b111101000;assign rom[9055] = 'b101001111;assign rom[9056] = 'b000111010;assign rom[9057] = 'b101110110;assign rom[9058] = 'b101100010;assign rom[9059] = 'b101001100;assign rom[9060] = 'b001001010;assign rom[9061] = 'b111011010;assign rom[9062] = 'b111011010;assign rom[9063] = 'b111011010;assign rom[9064] = 'b111011010;assign rom[9065] = 'b111011000;assign rom[9066] = 'b111011000;assign rom[9067] = 'b111011000;assign rom[9068] = 'b111011000;assign rom[9069] = 'b101111000;assign rom[9070] = 'b000110011;assign rom[9071] = 'b110000010;assign rom[9072] = 'b001101010;assign rom[9073] = 'b001011000;assign rom[9074] = 'b101001000;assign rom[9075] = 'b000101011;assign rom[9076] = 'b110000010;assign rom[9077] = 'b111000000;assign rom[9078] = 'b101001100;assign rom[9079] = 'b001001010;assign rom[9080] = 'b111111000;assign rom[9081] = 'b111101000;assign rom[9082] = 'b101001111;assign rom[9083] = 'b000111010;assign rom[9084] = 'b101110110;assign rom[9085] = 'b101100010;assign rom[9086] = 'b101001100;assign rom[9087] = 'b001001010;assign rom[9088] = 'b111011010;assign rom[9089] = 'b111011010;assign rom[9090] = 'b111011010;assign rom[9091] = 'b111011010;assign rom[9092] = 'b111011000;assign rom[9093] = 'b111011000;assign rom[9094] = 'b111011000;assign rom[9095] = 'b111011000;assign rom[9096] = 'b101111000;assign rom[9097] = 'b000110011;assign rom[9098] = 'b110000010;assign rom[9099] = 'b001101010;assign rom[9100] = 'b001011000;assign rom[9101] = 'b101001000;assign rom[9102] = 'b000101011;assign rom[9103] = 'b110000010;assign rom[9104] = 'b111000000;assign rom[9105] = 'b101001100;assign rom[9106] = 'b001001010;assign rom[9107] = 'b111111000;assign rom[9108] = 'b111101000;assign rom[9109] = 'b101001111;assign rom[9110] = 'b000111010;assign rom[9111] = 'b101110110;assign rom[9112] = 'b101100010;assign rom[9113] = 'b101001100;assign rom[9114] = 'b001001010;assign rom[9115] = 'b111011010;assign rom[9116] = 'b111011010;assign rom[9117] = 'b111011010;assign rom[9118] = 'b111011010;assign rom[9119] = 'b111011000;assign rom[9120] = 'b111011000;assign rom[9121] = 'b111011000;assign rom[9122] = 'b111011000;assign rom[9123] = 'b101111000;assign rom[9124] = 'b000110011;assign rom[9125] = 'b110000010;assign rom[9126] = 'b001101010;assign rom[9127] = 'b001011000;assign rom[9128] = 'b101001000;assign rom[9129] = 'b000101011;assign rom[9130] = 'b110000010;assign rom[9131] = 'b111000000;assign rom[9132] = 'b101001100;assign rom[9133] = 'b001001010;assign rom[9134] = 'b111111000;assign rom[9135] = 'b111101000;assign rom[9136] = 'b101001111;assign rom[9137] = 'b000111010;assign rom[9138] = 'b101110110;assign rom[9139] = 'b101100010;assign rom[9140] = 'b101001100;assign rom[9141] = 'b001001010;assign rom[9142] = 'b111011010;assign rom[9143] = 'b111011010;assign rom[9144] = 'b111011010;assign rom[9145] = 'b111011010;assign rom[9146] = 'b111011000;assign rom[9147] = 'b111011000;assign rom[9148] = 'b111011000;assign rom[9149] = 'b111011000;assign rom[9150] = 'b101111000;assign rom[9151] = 'b000110011;assign rom[9152] = 'b110000010;assign rom[9153] = 'b001101010;assign rom[9154] = 'b001011000;assign rom[9155] = 'b101001000;assign rom[9156] = 'b000101011;assign rom[9157] = 'b110000010;assign rom[9158] = 'b111000000;assign rom[9159] = 'b101001100;assign rom[9160] = 'b001001010;assign rom[9161] = 'b001000110;assign rom[9162] = 'b001100100;assign rom[9163] = 'b101100010;assign rom[9164] = 'b101001100;assign rom[9165] = 'b001001010;assign rom[9166] = 'b111011010;assign rom[9167] = 'b111011010;assign rom[9168] = 'b111011010;assign rom[9169] = 'b111011010;assign rom[9170] = 'b111011000;assign rom[9171] = 'b111011000;assign rom[9172] = 'b111011000;assign rom[9173] = 'b111011000;assign rom[9174] = 'b101111000;assign rom[9175] = 'b000110011;assign rom[9176] = 'b110000010;assign rom[9177] = 'b001101010;assign rom[9178] = 'b001011000;assign rom[9179] = 'b101001000;assign rom[9180] = 'b000101011;assign rom[9181] = 'b110000010;assign rom[9182] = 'b111000000;assign rom[9183] = 'b101001100;assign rom[9184] = 'b001001010;assign rom[9185] = 'b111111000;assign rom[9186] = 'b111101000;assign rom[9187] = 'b101001111;assign rom[9188] = 'b000111010;assign rom[9189] = 'b101110110;assign rom[9190] = 'b101100010;assign rom[9191] = 'b101001100;assign rom[9192] = 'b001001010;assign rom[9193] = 'b111011010;assign rom[9194] = 'b111011010;assign rom[9195] = 'b111011010;assign rom[9196] = 'b111011010;assign rom[9197] = 'b111011000;assign rom[9198] = 'b111011000;assign rom[9199] = 'b111011000;assign rom[9200] = 'b111011000;assign rom[9201] = 'b101111000;assign rom[9202] = 'b000110011;assign rom[9203] = 'b110000010;assign rom[9204] = 'b001101010;assign rom[9205] = 'b001011000;assign rom[9206] = 'b101001000;assign rom[9207] = 'b000101011;assign rom[9208] = 'b110000010;assign rom[9209] = 'b111000000;assign rom[9210] = 'b101001100;assign rom[9211] = 'b001001010;assign rom[9212] = 'b111111000;assign rom[9213] = 'b111101000;assign rom[9214] = 'b101001111;assign rom[9215] = 'b000111010;assign rom[9216] = 'b101110110;assign rom[9217] = 'b101100010;assign rom[9218] = 'b101001100;assign rom[9219] = 'b001001010;assign rom[9220] = 'b111011010;assign rom[9221] = 'b111011010;assign rom[9222] = 'b111011010;assign rom[9223] = 'b111011010;assign rom[9224] = 'b111011000;assign rom[9225] = 'b111011000;assign rom[9226] = 'b111011000;assign rom[9227] = 'b111011000;assign rom[9228] = 'b101111000;assign rom[9229] = 'b000110011;assign rom[9230] = 'b110000010;assign rom[9231] = 'b001101010;assign rom[9232] = 'b001011000;assign rom[9233] = 'b101001000;assign rom[9234] = 'b000101011;assign rom[9235] = 'b110000010;assign rom[9236] = 'b111000000;assign rom[9237] = 'b101001100;assign rom[9238] = 'b001001010;assign rom[9239] = 'b111111000;assign rom[9240] = 'b111101000;assign rom[9241] = 'b101001111;assign rom[9242] = 'b000111010;assign rom[9243] = 'b101110110;assign rom[9244] = 'b101100010;assign rom[9245] = 'b101001100;assign rom[9246] = 'b001001010;assign rom[9247] = 'b111011010;assign rom[9248] = 'b111011010;assign rom[9249] = 'b111011010;assign rom[9250] = 'b111011010;assign rom[9251] = 'b111011000;assign rom[9252] = 'b111011000;assign rom[9253] = 'b111011000;assign rom[9254] = 'b111011000;assign rom[9255] = 'b101111000;assign rom[9256] = 'b000110011;assign rom[9257] = 'b110000010;assign rom[9258] = 'b001101010;assign rom[9259] = 'b001011000;assign rom[9260] = 'b101001000;assign rom[9261] = 'b000101011;assign rom[9262] = 'b110000010;assign rom[9263] = 'b111000000;assign rom[9264] = 'b101001100;assign rom[9265] = 'b001001010;assign rom[9266] = 'b111111000;assign rom[9267] = 'b111101000;assign rom[9268] = 'b101001111;assign rom[9269] = 'b000111010;assign rom[9270] = 'b101110110;assign rom[9271] = 'b101100010;assign rom[9272] = 'b101001100;assign rom[9273] = 'b001001010;assign rom[9274] = 'b111011010;assign rom[9275] = 'b111011010;assign rom[9276] = 'b111011010;assign rom[9277] = 'b111011010;assign rom[9278] = 'b111011000;assign rom[9279] = 'b111011000;assign rom[9280] = 'b111011000;assign rom[9281] = 'b111011000;assign rom[9282] = 'b101111000;assign rom[9283] = 'b000110011;assign rom[9284] = 'b110000010;assign rom[9285] = 'b001101010;assign rom[9286] = 'b001011000;assign rom[9287] = 'b101001000;assign rom[9288] = 'b000101011;assign rom[9289] = 'b110000010;assign rom[9290] = 'b111000000;assign rom[9291] = 'b101001100;assign rom[9292] = 'b001001010;assign rom[9293] = 'b111111000;assign rom[9294] = 'b111101000;assign rom[9295] = 'b101001111;assign rom[9296] = 'b000111010;assign rom[9297] = 'b101110110;assign rom[9298] = 'b101100010;assign rom[9299] = 'b101001100;assign rom[9300] = 'b001001010;assign rom[9301] = 'b111011010;assign rom[9302] = 'b111011010;assign rom[9303] = 'b111011010;assign rom[9304] = 'b111011010;assign rom[9305] = 'b111011000;assign rom[9306] = 'b111011000;assign rom[9307] = 'b111011000;assign rom[9308] = 'b111011000;assign rom[9309] = 'b101111000;assign rom[9310] = 'b000110011;assign rom[9311] = 'b110000010;assign rom[9312] = 'b001101010;assign rom[9313] = 'b001011000;assign rom[9314] = 'b101001000;assign rom[9315] = 'b000101011;assign rom[9316] = 'b110000010;assign rom[9317] = 'b111000000;assign rom[9318] = 'b101001100;assign rom[9319] = 'b001001010;assign rom[9320] = 'b111111000;assign rom[9321] = 'b111101000;assign rom[9322] = 'b101001111;assign rom[9323] = 'b000111010;assign rom[9324] = 'b101110110;assign rom[9325] = 'b101100010;assign rom[9326] = 'b101001100;assign rom[9327] = 'b001001010;assign rom[9328] = 'b111011010;assign rom[9329] = 'b111011010;assign rom[9330] = 'b111011010;assign rom[9331] = 'b111011010;assign rom[9332] = 'b111011000;assign rom[9333] = 'b111011000;assign rom[9334] = 'b111011000;assign rom[9335] = 'b111011000;assign rom[9336] = 'b101111000;assign rom[9337] = 'b000110011;assign rom[9338] = 'b110000010;assign rom[9339] = 'b001101010;assign rom[9340] = 'b001011000;assign rom[9341] = 'b101001000;assign rom[9342] = 'b000101011;assign rom[9343] = 'b110000010;assign rom[9344] = 'b111000000;assign rom[9345] = 'b101001100;assign rom[9346] = 'b001001010;assign rom[9347] = 'b111111000;assign rom[9348] = 'b111101000;assign rom[9349] = 'b101001111;assign rom[9350] = 'b000111010;assign rom[9351] = 'b101110110;assign rom[9352] = 'b101100010;assign rom[9353] = 'b101001100;assign rom[9354] = 'b001001010;assign rom[9355] = 'b111011010;assign rom[9356] = 'b111011010;assign rom[9357] = 'b111011010;assign rom[9358] = 'b111011010;assign rom[9359] = 'b111011000;assign rom[9360] = 'b111011000;assign rom[9361] = 'b111011000;assign rom[9362] = 'b111011000;assign rom[9363] = 'b101111000;assign rom[9364] = 'b000110011;assign rom[9365] = 'b110000010;assign rom[9366] = 'b001101010;assign rom[9367] = 'b001011000;assign rom[9368] = 'b101001000;assign rom[9369] = 'b000101011;assign rom[9370] = 'b110000010;assign rom[9371] = 'b111000000;assign rom[9372] = 'b101001100;assign rom[9373] = 'b001001010;assign rom[9374] = 'b111111000;assign rom[9375] = 'b111101000;assign rom[9376] = 'b101001111;assign rom[9377] = 'b000111010;assign rom[9378] = 'b101110110;assign rom[9379] = 'b101100010;assign rom[9380] = 'b101001100;assign rom[9381] = 'b001001010;assign rom[9382] = 'b111011010;assign rom[9383] = 'b111011010;assign rom[9384] = 'b111011010;assign rom[9385] = 'b111011010;assign rom[9386] = 'b111011000;assign rom[9387] = 'b111011000;assign rom[9388] = 'b111011000;assign rom[9389] = 'b111011000;assign rom[9390] = 'b101111000;assign rom[9391] = 'b000110011;assign rom[9392] = 'b110000010;assign rom[9393] = 'b001101010;assign rom[9394] = 'b001011000;assign rom[9395] = 'b101001000;assign rom[9396] = 'b000101011;assign rom[9397] = 'b110000010;assign rom[9398] = 'b111000000;assign rom[9399] = 'b101001100;assign rom[9400] = 'b001001010;assign rom[9401] = 'b001000110;assign rom[9402] = 'b001100100;assign rom[9403] = 'b101100010;assign rom[9404] = 'b101001100;assign rom[9405] = 'b001001010;assign rom[9406] = 'b111011010;assign rom[9407] = 'b111011010;assign rom[9408] = 'b111011010;assign rom[9409] = 'b111011010;assign rom[9410] = 'b111011000;assign rom[9411] = 'b111011000;assign rom[9412] = 'b111011000;assign rom[9413] = 'b111011000;assign rom[9414] = 'b101111000;assign rom[9415] = 'b000110011;assign rom[9416] = 'b110000010;assign rom[9417] = 'b001101010;assign rom[9418] = 'b001011000;assign rom[9419] = 'b101001000;assign rom[9420] = 'b000101011;assign rom[9421] = 'b110000010;assign rom[9422] = 'b111000000;assign rom[9423] = 'b101001100;assign rom[9424] = 'b001001010;assign rom[9425] = 'b111111000;assign rom[9426] = 'b111101000;assign rom[9427] = 'b101001111;assign rom[9428] = 'b000111010;assign rom[9429] = 'b101110110;assign rom[9430] = 'b101100010;assign rom[9431] = 'b101001100;assign rom[9432] = 'b001001010;assign rom[9433] = 'b111011010;assign rom[9434] = 'b111011010;assign rom[9435] = 'b111011010;assign rom[9436] = 'b111011010;assign rom[9437] = 'b111011000;assign rom[9438] = 'b111011000;assign rom[9439] = 'b111011000;assign rom[9440] = 'b111011000;assign rom[9441] = 'b101111000;assign rom[9442] = 'b000110011;assign rom[9443] = 'b110000010;assign rom[9444] = 'b001101010;assign rom[9445] = 'b001011000;assign rom[9446] = 'b101001000;assign rom[9447] = 'b000101011;assign rom[9448] = 'b110000010;assign rom[9449] = 'b111000000;assign rom[9450] = 'b101001100;assign rom[9451] = 'b001001010;assign rom[9452] = 'b111111000;assign rom[9453] = 'b111101000;assign rom[9454] = 'b101001111;assign rom[9455] = 'b000111010;assign rom[9456] = 'b101110110;assign rom[9457] = 'b101100010;assign rom[9458] = 'b101001100;assign rom[9459] = 'b001001010;assign rom[9460] = 'b111011010;assign rom[9461] = 'b111011010;assign rom[9462] = 'b111011010;assign rom[9463] = 'b111011010;assign rom[9464] = 'b111011000;assign rom[9465] = 'b111011000;assign rom[9466] = 'b111011000;assign rom[9467] = 'b111011000;assign rom[9468] = 'b101111000;assign rom[9469] = 'b000110011;assign rom[9470] = 'b110000010;assign rom[9471] = 'b001101010;assign rom[9472] = 'b001011000;assign rom[9473] = 'b101001000;assign rom[9474] = 'b000101011;assign rom[9475] = 'b110000010;assign rom[9476] = 'b111000000;assign rom[9477] = 'b101001100;assign rom[9478] = 'b001001010;assign rom[9479] = 'b111111000;assign rom[9480] = 'b111101000;assign rom[9481] = 'b101001111;assign rom[9482] = 'b000111010;assign rom[9483] = 'b101110110;assign rom[9484] = 'b101100010;assign rom[9485] = 'b101001100;assign rom[9486] = 'b001001010;assign rom[9487] = 'b111011010;assign rom[9488] = 'b111011010;assign rom[9489] = 'b111011010;assign rom[9490] = 'b111011010;assign rom[9491] = 'b111011000;assign rom[9492] = 'b111011000;assign rom[9493] = 'b111011000;assign rom[9494] = 'b111011000;assign rom[9495] = 'b101111000;assign rom[9496] = 'b000110011;assign rom[9497] = 'b110000010;assign rom[9498] = 'b001101010;assign rom[9499] = 'b001011000;assign rom[9500] = 'b101001000;assign rom[9501] = 'b000101011;assign rom[9502] = 'b110000010;assign rom[9503] = 'b111000000;assign rom[9504] = 'b101001100;assign rom[9505] = 'b001001010;assign rom[9506] = 'b111111000;assign rom[9507] = 'b111101000;assign rom[9508] = 'b101001111;assign rom[9509] = 'b000111010;assign rom[9510] = 'b101110110;assign rom[9511] = 'b101100010;assign rom[9512] = 'b101001100;assign rom[9513] = 'b001001010;assign rom[9514] = 'b111011010;assign rom[9515] = 'b111011010;assign rom[9516] = 'b111011010;assign rom[9517] = 'b111011010;assign rom[9518] = 'b111011000;assign rom[9519] = 'b111011000;assign rom[9520] = 'b111011000;assign rom[9521] = 'b111011000;assign rom[9522] = 'b101111000;assign rom[9523] = 'b000110011;assign rom[9524] = 'b110000010;assign rom[9525] = 'b001101010;assign rom[9526] = 'b001011000;assign rom[9527] = 'b101001000;assign rom[9528] = 'b000101011;assign rom[9529] = 'b110000010;assign rom[9530] = 'b111000000;assign rom[9531] = 'b101001100;assign rom[9532] = 'b001001010;assign rom[9533] = 'b111111000;assign rom[9534] = 'b111101000;assign rom[9535] = 'b101001111;assign rom[9536] = 'b000111010;assign rom[9537] = 'b101110110;assign rom[9538] = 'b101100010;assign rom[9539] = 'b101001100;assign rom[9540] = 'b001001010;assign rom[9541] = 'b111011010;assign rom[9542] = 'b111011010;assign rom[9543] = 'b111011010;assign rom[9544] = 'b111011010;assign rom[9545] = 'b111011000;assign rom[9546] = 'b111011000;assign rom[9547] = 'b111011000;assign rom[9548] = 'b111011000;assign rom[9549] = 'b101111000;assign rom[9550] = 'b000110011;assign rom[9551] = 'b110000010;assign rom[9552] = 'b001101010;assign rom[9553] = 'b001011000;assign rom[9554] = 'b101001000;assign rom[9555] = 'b000101011;assign rom[9556] = 'b110000010;assign rom[9557] = 'b111000000;assign rom[9558] = 'b101001100;assign rom[9559] = 'b001001010;assign rom[9560] = 'b111111000;assign rom[9561] = 'b111101000;assign rom[9562] = 'b101001111;assign rom[9563] = 'b000111010;assign rom[9564] = 'b101110110;assign rom[9565] = 'b101100010;assign rom[9566] = 'b101001100;assign rom[9567] = 'b001001010;assign rom[9568] = 'b111011010;assign rom[9569] = 'b111011010;assign rom[9570] = 'b111011010;assign rom[9571] = 'b111011010;assign rom[9572] = 'b111011000;assign rom[9573] = 'b111011000;assign rom[9574] = 'b111011000;assign rom[9575] = 'b111011000;assign rom[9576] = 'b101111000;assign rom[9577] = 'b000110011;assign rom[9578] = 'b110000010;assign rom[9579] = 'b001101010;assign rom[9580] = 'b001011000;assign rom[9581] = 'b101001000;assign rom[9582] = 'b000101011;assign rom[9583] = 'b110000010;assign rom[9584] = 'b111000000;assign rom[9585] = 'b101001100;assign rom[9586] = 'b001001010;assign rom[9587] = 'b111111000;assign rom[9588] = 'b111101000;assign rom[9589] = 'b101001111;assign rom[9590] = 'b000111010;assign rom[9591] = 'b101110110;assign rom[9592] = 'b101100010;assign rom[9593] = 'b101001100;assign rom[9594] = 'b001001010;assign rom[9595] = 'b111011010;assign rom[9596] = 'b111011010;assign rom[9597] = 'b111011010;assign rom[9598] = 'b111011010;assign rom[9599] = 'b111011000;assign rom[9600] = 'b111011000;assign rom[9601] = 'b111011000;assign rom[9602] = 'b111011000;assign rom[9603] = 'b101111000;assign rom[9604] = 'b000110011;assign rom[9605] = 'b110000010;assign rom[9606] = 'b001101010;assign rom[9607] = 'b001011000;assign rom[9608] = 'b101001000;assign rom[9609] = 'b000101011;assign rom[9610] = 'b110000010;assign rom[9611] = 'b111000000;assign rom[9612] = 'b101001100;assign rom[9613] = 'b001001010;assign rom[9614] = 'b111111000;assign rom[9615] = 'b111101000;assign rom[9616] = 'b101001111;assign rom[9617] = 'b000111010;assign rom[9618] = 'b101110110;assign rom[9619] = 'b101100010;assign rom[9620] = 'b101001100;assign rom[9621] = 'b001001010;assign rom[9622] = 'b111011010;assign rom[9623] = 'b111011010;assign rom[9624] = 'b111011010;assign rom[9625] = 'b111011010;assign rom[9626] = 'b111011000;assign rom[9627] = 'b111011000;assign rom[9628] = 'b111011000;assign rom[9629] = 'b111011000;assign rom[9630] = 'b101111000;assign rom[9631] = 'b000110011;assign rom[9632] = 'b110000010;assign rom[9633] = 'b001101010;assign rom[9634] = 'b001011000;assign rom[9635] = 'b101001000;assign rom[9636] = 'b000101011;assign rom[9637] = 'b110000010;assign rom[9638] = 'b111000000;assign rom[9639] = 'b101001100;assign rom[9640] = 'b001001010;assign rom[9641] = 'b001000110;assign rom[9642] = 'b001100100;assign rom[9643] = 'b101100010;assign rom[9644] = 'b101001100;assign rom[9645] = 'b001001010;assign rom[9646] = 'b111011010;assign rom[9647] = 'b111011010;assign rom[9648] = 'b111011010;assign rom[9649] = 'b111011010;assign rom[9650] = 'b111011000;assign rom[9651] = 'b111011000;assign rom[9652] = 'b111011000;assign rom[9653] = 'b111011000;assign rom[9654] = 'b101111000;assign rom[9655] = 'b000110011;assign rom[9656] = 'b110000010;assign rom[9657] = 'b001101010;assign rom[9658] = 'b001011000;assign rom[9659] = 'b101001000;assign rom[9660] = 'b000101011;assign rom[9661] = 'b110000010;assign rom[9662] = 'b111000000;assign rom[9663] = 'b101001100;assign rom[9664] = 'b001001010;assign rom[9665] = 'b111111000;assign rom[9666] = 'b111101000;assign rom[9667] = 'b101001111;assign rom[9668] = 'b000111010;assign rom[9669] = 'b101110110;assign rom[9670] = 'b101100010;assign rom[9671] = 'b101001100;assign rom[9672] = 'b001001010;assign rom[9673] = 'b111011010;assign rom[9674] = 'b111011010;assign rom[9675] = 'b111011010;assign rom[9676] = 'b111011010;assign rom[9677] = 'b111011000;assign rom[9678] = 'b111011000;assign rom[9679] = 'b111011000;assign rom[9680] = 'b111011000;assign rom[9681] = 'b101111000;assign rom[9682] = 'b000110011;assign rom[9683] = 'b110000010;assign rom[9684] = 'b001101010;assign rom[9685] = 'b001011000;assign rom[9686] = 'b101001000;assign rom[9687] = 'b000101011;assign rom[9688] = 'b110000010;assign rom[9689] = 'b111000000;assign rom[9690] = 'b101001100;assign rom[9691] = 'b001001010;assign rom[9692] = 'b111111000;assign rom[9693] = 'b111101000;assign rom[9694] = 'b101001111;assign rom[9695] = 'b000111010;assign rom[9696] = 'b101110110;assign rom[9697] = 'b101100010;assign rom[9698] = 'b101001100;assign rom[9699] = 'b001001010;assign rom[9700] = 'b111011010;assign rom[9701] = 'b111011010;assign rom[9702] = 'b111011010;assign rom[9703] = 'b111011010;assign rom[9704] = 'b111011000;assign rom[9705] = 'b111011000;assign rom[9706] = 'b111011000;assign rom[9707] = 'b111011000;assign rom[9708] = 'b101111000;assign rom[9709] = 'b000110011;assign rom[9710] = 'b110000010;assign rom[9711] = 'b001101010;assign rom[9712] = 'b001011000;assign rom[9713] = 'b101001000;assign rom[9714] = 'b000101011;assign rom[9715] = 'b110000010;assign rom[9716] = 'b111000000;assign rom[9717] = 'b101001100;assign rom[9718] = 'b001001010;assign rom[9719] = 'b111111000;assign rom[9720] = 'b111101000;assign rom[9721] = 'b101001111;assign rom[9722] = 'b000111010;assign rom[9723] = 'b101110110;assign rom[9724] = 'b101100010;assign rom[9725] = 'b101001100;assign rom[9726] = 'b001001010;assign rom[9727] = 'b111011010;assign rom[9728] = 'b111011010;assign rom[9729] = 'b111011010;assign rom[9730] = 'b111011010;assign rom[9731] = 'b111011000;assign rom[9732] = 'b111011000;assign rom[9733] = 'b111011000;assign rom[9734] = 'b111011000;assign rom[9735] = 'b101111000;assign rom[9736] = 'b000110011;assign rom[9737] = 'b110000010;assign rom[9738] = 'b001101010;assign rom[9739] = 'b001011000;assign rom[9740] = 'b101001000;assign rom[9741] = 'b000101011;assign rom[9742] = 'b110000010;assign rom[9743] = 'b111000000;assign rom[9744] = 'b101001100;assign rom[9745] = 'b001001010;assign rom[9746] = 'b111111000;assign rom[9747] = 'b111101000;assign rom[9748] = 'b101001111;assign rom[9749] = 'b000111010;assign rom[9750] = 'b101110110;assign rom[9751] = 'b101100010;assign rom[9752] = 'b101001100;assign rom[9753] = 'b001001010;assign rom[9754] = 'b111011010;assign rom[9755] = 'b111011010;assign rom[9756] = 'b111011010;assign rom[9757] = 'b111011010;assign rom[9758] = 'b111011000;assign rom[9759] = 'b111011000;assign rom[9760] = 'b111011000;assign rom[9761] = 'b111011000;assign rom[9762] = 'b101111000;assign rom[9763] = 'b000110011;assign rom[9764] = 'b110000010;assign rom[9765] = 'b001101010;assign rom[9766] = 'b001011000;assign rom[9767] = 'b101001000;assign rom[9768] = 'b000101011;assign rom[9769] = 'b110000010;assign rom[9770] = 'b111000000;assign rom[9771] = 'b101001100;assign rom[9772] = 'b001001010;assign rom[9773] = 'b111111000;assign rom[9774] = 'b111101000;assign rom[9775] = 'b101001111;assign rom[9776] = 'b000111010;assign rom[9777] = 'b101110110;assign rom[9778] = 'b101100010;assign rom[9779] = 'b101001100;assign rom[9780] = 'b001001010;assign rom[9781] = 'b111011010;assign rom[9782] = 'b111011010;assign rom[9783] = 'b111011010;assign rom[9784] = 'b111011010;assign rom[9785] = 'b111011000;assign rom[9786] = 'b111011000;assign rom[9787] = 'b111011000;assign rom[9788] = 'b111011000;assign rom[9789] = 'b101111000;assign rom[9790] = 'b000110011;assign rom[9791] = 'b110000010;assign rom[9792] = 'b001101010;assign rom[9793] = 'b001011000;assign rom[9794] = 'b101001000;assign rom[9795] = 'b000101011;assign rom[9796] = 'b110000010;assign rom[9797] = 'b111000000;assign rom[9798] = 'b101001100;assign rom[9799] = 'b001001010;assign rom[9800] = 'b111111000;assign rom[9801] = 'b111101000;assign rom[9802] = 'b101001111;assign rom[9803] = 'b000111010;assign rom[9804] = 'b101110110;assign rom[9805] = 'b101100010;assign rom[9806] = 'b101001100;assign rom[9807] = 'b001001010;assign rom[9808] = 'b111011010;assign rom[9809] = 'b111011010;assign rom[9810] = 'b111011010;assign rom[9811] = 'b111011010;assign rom[9812] = 'b111011000;assign rom[9813] = 'b111011000;assign rom[9814] = 'b111011000;assign rom[9815] = 'b111011000;assign rom[9816] = 'b101111000;assign rom[9817] = 'b000110011;assign rom[9818] = 'b110000010;assign rom[9819] = 'b001101010;assign rom[9820] = 'b001011000;assign rom[9821] = 'b101001000;assign rom[9822] = 'b000101011;assign rom[9823] = 'b110000010;assign rom[9824] = 'b111000000;assign rom[9825] = 'b101001100;assign rom[9826] = 'b001001010;assign rom[9827] = 'b111111000;assign rom[9828] = 'b111101000;assign rom[9829] = 'b101001111;assign rom[9830] = 'b000111010;assign rom[9831] = 'b101110110;assign rom[9832] = 'b101100010;assign rom[9833] = 'b101001100;assign rom[9834] = 'b001001010;assign rom[9835] = 'b111011010;assign rom[9836] = 'b111011010;assign rom[9837] = 'b111011010;assign rom[9838] = 'b111011010;assign rom[9839] = 'b111011000;assign rom[9840] = 'b111011000;assign rom[9841] = 'b111011000;assign rom[9842] = 'b111011000;assign rom[9843] = 'b101111000;assign rom[9844] = 'b000110011;assign rom[9845] = 'b110000010;assign rom[9846] = 'b001101010;assign rom[9847] = 'b001011000;assign rom[9848] = 'b101001000;assign rom[9849] = 'b000101011;assign rom[9850] = 'b110000010;assign rom[9851] = 'b111000000;assign rom[9852] = 'b101001100;assign rom[9853] = 'b001001010;assign rom[9854] = 'b111111000;assign rom[9855] = 'b111101000;assign rom[9856] = 'b101001111;assign rom[9857] = 'b000111010;assign rom[9858] = 'b101110110;assign rom[9859] = 'b101100010;assign rom[9860] = 'b101001100;assign rom[9861] = 'b001001010;assign rom[9862] = 'b111011010;assign rom[9863] = 'b111011010;assign rom[9864] = 'b111011010;assign rom[9865] = 'b111011010;assign rom[9866] = 'b111011000;assign rom[9867] = 'b111011000;assign rom[9868] = 'b111011000;assign rom[9869] = 'b111011000;assign rom[9870] = 'b101111000;assign rom[9871] = 'b000110011;assign rom[9872] = 'b110000010;assign rom[9873] = 'b001101010;assign rom[9874] = 'b001011000;assign rom[9875] = 'b101001000;assign rom[9876] = 'b000101011;assign rom[9877] = 'b110000010;assign rom[9878] = 'b111000000;assign rom[9879] = 'b101001100;assign rom[9880] = 'b001001010;assign rom[9881] = 'b001000110;assign rom[9882] = 'b001100100;assign rom[9883] = 'b101100010;assign rom[9884] = 'b101001100;assign rom[9885] = 'b001001010;assign rom[9886] = 'b111011010;assign rom[9887] = 'b111011010;assign rom[9888] = 'b111011010;assign rom[9889] = 'b111011010;assign rom[9890] = 'b111011000;assign rom[9891] = 'b111011000;assign rom[9892] = 'b111011000;assign rom[9893] = 'b111011000;assign rom[9894] = 'b101111000;assign rom[9895] = 'b000110011;assign rom[9896] = 'b110000010;assign rom[9897] = 'b001101010;assign rom[9898] = 'b001011000;assign rom[9899] = 'b101001000;assign rom[9900] = 'b000101011;assign rom[9901] = 'b110000010;assign rom[9902] = 'b111000000;assign rom[9903] = 'b101001100;assign rom[9904] = 'b001001010;assign rom[9905] = 'b111111000;assign rom[9906] = 'b111101000;assign rom[9907] = 'b101001111;assign rom[9908] = 'b000111010;assign rom[9909] = 'b101110110;assign rom[9910] = 'b101100010;assign rom[9911] = 'b101001100;assign rom[9912] = 'b001001010;assign rom[9913] = 'b111011010;assign rom[9914] = 'b111011010;assign rom[9915] = 'b111011010;assign rom[9916] = 'b111011010;assign rom[9917] = 'b111011000;assign rom[9918] = 'b111011000;assign rom[9919] = 'b111011000;assign rom[9920] = 'b111011000;assign rom[9921] = 'b101111000;assign rom[9922] = 'b000110011;assign rom[9923] = 'b110000010;assign rom[9924] = 'b001101010;assign rom[9925] = 'b001011000;assign rom[9926] = 'b101001000;assign rom[9927] = 'b000101011;assign rom[9928] = 'b110000010;assign rom[9929] = 'b111000000;assign rom[9930] = 'b101001100;assign rom[9931] = 'b001001010;assign rom[9932] = 'b111111000;assign rom[9933] = 'b111101000;assign rom[9934] = 'b101001111;assign rom[9935] = 'b000111010;assign rom[9936] = 'b101110110;assign rom[9937] = 'b101100010;assign rom[9938] = 'b101001100;assign rom[9939] = 'b001001010;assign rom[9940] = 'b111011010;assign rom[9941] = 'b111011010;assign rom[9942] = 'b111011010;assign rom[9943] = 'b111011010;assign rom[9944] = 'b111011000;assign rom[9945] = 'b111011000;assign rom[9946] = 'b111011000;assign rom[9947] = 'b111011000;assign rom[9948] = 'b101111000;assign rom[9949] = 'b000110011;assign rom[9950] = 'b110000010;assign rom[9951] = 'b001101010;assign rom[9952] = 'b001011000;assign rom[9953] = 'b101001000;assign rom[9954] = 'b000101011;assign rom[9955] = 'b110000010;assign rom[9956] = 'b111000000;assign rom[9957] = 'b101001100;assign rom[9958] = 'b001001010;assign rom[9959] = 'b111111000;assign rom[9960] = 'b111101000;assign rom[9961] = 'b101001111;assign rom[9962] = 'b000111010;assign rom[9963] = 'b101110110;assign rom[9964] = 'b101100010;assign rom[9965] = 'b101001100;assign rom[9966] = 'b001001010;assign rom[9967] = 'b111011010;assign rom[9968] = 'b111011010;assign rom[9969] = 'b111011010;assign rom[9970] = 'b111011010;assign rom[9971] = 'b111011000;assign rom[9972] = 'b111011000;assign rom[9973] = 'b111011000;assign rom[9974] = 'b111011000;assign rom[9975] = 'b101111000;assign rom[9976] = 'b000110011;assign rom[9977] = 'b110000010;assign rom[9978] = 'b001101010;assign rom[9979] = 'b001011000;assign rom[9980] = 'b101001000;assign rom[9981] = 'b000101011;assign rom[9982] = 'b110000010;assign rom[9983] = 'b111000000;assign rom[9984] = 'b101001100;assign rom[9985] = 'b001001010;assign rom[9986] = 'b111111000;assign rom[9987] = 'b111101000;assign rom[9988] = 'b101001111;assign rom[9989] = 'b000111010;assign rom[9990] = 'b101110110;assign rom[9991] = 'b101100010;assign rom[9992] = 'b101001100;assign rom[9993] = 'b001001010;assign rom[9994] = 'b111011010;assign rom[9995] = 'b111011010;assign rom[9996] = 'b111011010;assign rom[9997] = 'b111011010;assign rom[9998] = 'b111011000;assign rom[9999] = 'b111011000;assign rom[10000] = 'b111011000;assign rom[10001] = 'b111011000;assign rom[10002] = 'b101111000;assign rom[10003] = 'b000110011;assign rom[10004] = 'b110000010;assign rom[10005] = 'b001101010;assign rom[10006] = 'b001011000;assign rom[10007] = 'b101001000;assign rom[10008] = 'b000101011;assign rom[10009] = 'b110000010;assign rom[10010] = 'b111000000;assign rom[10011] = 'b101001100;assign rom[10012] = 'b001001010;assign rom[10013] = 'b111111000;assign rom[10014] = 'b111101000;assign rom[10015] = 'b101001111;assign rom[10016] = 'b000111010;assign rom[10017] = 'b101110110;assign rom[10018] = 'b101100010;assign rom[10019] = 'b101001100;assign rom[10020] = 'b001001010;assign rom[10021] = 'b111011010;assign rom[10022] = 'b111011010;assign rom[10023] = 'b111011010;assign rom[10024] = 'b111011010;assign rom[10025] = 'b111011000;assign rom[10026] = 'b111011000;assign rom[10027] = 'b111011000;assign rom[10028] = 'b111011000;assign rom[10029] = 'b101111000;assign rom[10030] = 'b000110011;assign rom[10031] = 'b110000010;assign rom[10032] = 'b001101010;assign rom[10033] = 'b001011000;assign rom[10034] = 'b101001000;assign rom[10035] = 'b000101011;assign rom[10036] = 'b110000010;assign rom[10037] = 'b111000000;assign rom[10038] = 'b101001100;assign rom[10039] = 'b001001010;assign rom[10040] = 'b111111000;assign rom[10041] = 'b111101000;assign rom[10042] = 'b101001111;assign rom[10043] = 'b000111010;assign rom[10044] = 'b101110110;assign rom[10045] = 'b101100010;assign rom[10046] = 'b101001100;assign rom[10047] = 'b001001010;assign rom[10048] = 'b111011010;assign rom[10049] = 'b111011010;assign rom[10050] = 'b111011010;assign rom[10051] = 'b111011010;assign rom[10052] = 'b111011000;assign rom[10053] = 'b111011000;assign rom[10054] = 'b111011000;assign rom[10055] = 'b111011000;assign rom[10056] = 'b101111000;assign rom[10057] = 'b000110011;assign rom[10058] = 'b110000010;assign rom[10059] = 'b001101010;assign rom[10060] = 'b001011000;assign rom[10061] = 'b101001000;assign rom[10062] = 'b000101011;assign rom[10063] = 'b110000010;assign rom[10064] = 'b111000000;assign rom[10065] = 'b101001100;assign rom[10066] = 'b001001010;assign rom[10067] = 'b111111000;assign rom[10068] = 'b111101000;assign rom[10069] = 'b101001111;assign rom[10070] = 'b000111010;assign rom[10071] = 'b101110110;assign rom[10072] = 'b101100010;assign rom[10073] = 'b101001100;assign rom[10074] = 'b001001010;assign rom[10075] = 'b111011010;assign rom[10076] = 'b111011010;assign rom[10077] = 'b111011010;assign rom[10078] = 'b111011010;assign rom[10079] = 'b111011000;assign rom[10080] = 'b111011000;assign rom[10081] = 'b111011000;assign rom[10082] = 'b111011000;assign rom[10083] = 'b101111000;assign rom[10084] = 'b000110011;assign rom[10085] = 'b110000010;assign rom[10086] = 'b001101010;assign rom[10087] = 'b001011000;assign rom[10088] = 'b101001000;assign rom[10089] = 'b000101011;assign rom[10090] = 'b110000010;assign rom[10091] = 'b111000000;assign rom[10092] = 'b101001100;assign rom[10093] = 'b001001010;assign rom[10094] = 'b111111000;assign rom[10095] = 'b111101000;assign rom[10096] = 'b101001111;assign rom[10097] = 'b000111010;assign rom[10098] = 'b101110110;assign rom[10099] = 'b101100010;assign rom[10100] = 'b101001100;assign rom[10101] = 'b001001010;assign rom[10102] = 'b111011010;assign rom[10103] = 'b111011010;assign rom[10104] = 'b111011010;assign rom[10105] = 'b111011010;assign rom[10106] = 'b111011000;assign rom[10107] = 'b111011000;assign rom[10108] = 'b111011000;assign rom[10109] = 'b111011000;assign rom[10110] = 'b101111000;assign rom[10111] = 'b000110011;assign rom[10112] = 'b110000010;assign rom[10113] = 'b001101010;assign rom[10114] = 'b001011000;assign rom[10115] = 'b101001000;assign rom[10116] = 'b000101011;assign rom[10117] = 'b110000010;assign rom[10118] = 'b111000000;assign rom[10119] = 'b101001100;assign rom[10120] = 'b001001010;assign rom[10121] = 'b001000110;assign rom[10122] = 'b001100100;assign rom[10123] = 'b101100010;assign rom[10124] = 'b101001100;assign rom[10125] = 'b001001010;assign rom[10126] = 'b111011010;assign rom[10127] = 'b111011010;assign rom[10128] = 'b111011010;assign rom[10129] = 'b111011010;assign rom[10130] = 'b111011000;assign rom[10131] = 'b111011000;assign rom[10132] = 'b111011000;assign rom[10133] = 'b111011000;assign rom[10134] = 'b101111000;assign rom[10135] = 'b000110011;assign rom[10136] = 'b110000010;assign rom[10137] = 'b001101010;assign rom[10138] = 'b001011000;assign rom[10139] = 'b101001000;assign rom[10140] = 'b000101011;assign rom[10141] = 'b110000010;assign rom[10142] = 'b111000000;assign rom[10143] = 'b101001100;assign rom[10144] = 'b001001010;assign rom[10145] = 'b111111000;assign rom[10146] = 'b111101000;assign rom[10147] = 'b101001111;assign rom[10148] = 'b000111010;assign rom[10149] = 'b101110110;assign rom[10150] = 'b101100010;assign rom[10151] = 'b101001100;assign rom[10152] = 'b001001010;assign rom[10153] = 'b111011010;assign rom[10154] = 'b111011010;assign rom[10155] = 'b111011010;assign rom[10156] = 'b111011010;assign rom[10157] = 'b111011000;assign rom[10158] = 'b111011000;assign rom[10159] = 'b111011000;assign rom[10160] = 'b111011000;assign rom[10161] = 'b101111000;assign rom[10162] = 'b000110011;assign rom[10163] = 'b110000010;assign rom[10164] = 'b001101010;assign rom[10165] = 'b001011000;assign rom[10166] = 'b101001000;assign rom[10167] = 'b000101011;assign rom[10168] = 'b110000010;assign rom[10169] = 'b111000000;assign rom[10170] = 'b101001100;assign rom[10171] = 'b001001010;assign rom[10172] = 'b111111000;assign rom[10173] = 'b111101000;assign rom[10174] = 'b101001111;assign rom[10175] = 'b000111010;assign rom[10176] = 'b101110110;assign rom[10177] = 'b101100010;assign rom[10178] = 'b101001100;assign rom[10179] = 'b001001010;assign rom[10180] = 'b111011010;assign rom[10181] = 'b111011010;assign rom[10182] = 'b111011010;assign rom[10183] = 'b111011010;assign rom[10184] = 'b111011000;assign rom[10185] = 'b111011000;assign rom[10186] = 'b111011000;assign rom[10187] = 'b111011000;assign rom[10188] = 'b101111000;assign rom[10189] = 'b000110011;assign rom[10190] = 'b110000010;assign rom[10191] = 'b001101010;assign rom[10192] = 'b001011000;assign rom[10193] = 'b101001000;assign rom[10194] = 'b000101011;assign rom[10195] = 'b110000010;assign rom[10196] = 'b111000000;assign rom[10197] = 'b101001100;assign rom[10198] = 'b001001010;assign rom[10199] = 'b111111000;assign rom[10200] = 'b111101000;assign rom[10201] = 'b101001111;assign rom[10202] = 'b000111010;assign rom[10203] = 'b101110110;assign rom[10204] = 'b101100010;assign rom[10205] = 'b101001100;assign rom[10206] = 'b001001010;assign rom[10207] = 'b111011010;assign rom[10208] = 'b111011010;assign rom[10209] = 'b111011010;assign rom[10210] = 'b111011010;assign rom[10211] = 'b111011000;assign rom[10212] = 'b111011000;assign rom[10213] = 'b111011000;assign rom[10214] = 'b111011000;assign rom[10215] = 'b101111000;assign rom[10216] = 'b000110011;assign rom[10217] = 'b110000010;assign rom[10218] = 'b001101010;assign rom[10219] = 'b001011000;assign rom[10220] = 'b101001000;assign rom[10221] = 'b000101011;assign rom[10222] = 'b110000010;assign rom[10223] = 'b111000000;assign rom[10224] = 'b101001100;assign rom[10225] = 'b001001010;assign rom[10226] = 'b111111000;assign rom[10227] = 'b111101000;assign rom[10228] = 'b101001111;assign rom[10229] = 'b000111010;assign rom[10230] = 'b101110110;assign rom[10231] = 'b101100010;assign rom[10232] = 'b101001100;assign rom[10233] = 'b001001010;assign rom[10234] = 'b111011010;assign rom[10235] = 'b111011010;assign rom[10236] = 'b111011010;assign rom[10237] = 'b111011010;assign rom[10238] = 'b111011000;assign rom[10239] = 'b111011000;assign rom[10240] = 'b111011000;assign rom[10241] = 'b111011000;assign rom[10242] = 'b101111000;assign rom[10243] = 'b000110011;assign rom[10244] = 'b110000010;assign rom[10245] = 'b001101010;assign rom[10246] = 'b001011000;assign rom[10247] = 'b101001000;assign rom[10248] = 'b000101011;assign rom[10249] = 'b110000010;assign rom[10250] = 'b111000000;assign rom[10251] = 'b101001100;assign rom[10252] = 'b001001010;assign rom[10253] = 'b111111000;assign rom[10254] = 'b111101000;assign rom[10255] = 'b101001111;assign rom[10256] = 'b000111010;assign rom[10257] = 'b101110110;assign rom[10258] = 'b101100010;assign rom[10259] = 'b101001100;assign rom[10260] = 'b001001010;assign rom[10261] = 'b111011010;assign rom[10262] = 'b111011010;assign rom[10263] = 'b111011010;assign rom[10264] = 'b111011010;assign rom[10265] = 'b111011000;assign rom[10266] = 'b111011000;assign rom[10267] = 'b111011000;assign rom[10268] = 'b111011000;assign rom[10269] = 'b101111000;assign rom[10270] = 'b000110011;assign rom[10271] = 'b110000010;assign rom[10272] = 'b001101010;assign rom[10273] = 'b001011000;assign rom[10274] = 'b101001000;assign rom[10275] = 'b000101011;assign rom[10276] = 'b110000010;assign rom[10277] = 'b111000000;assign rom[10278] = 'b101001100;assign rom[10279] = 'b001001010;assign rom[10280] = 'b111111000;assign rom[10281] = 'b111101000;assign rom[10282] = 'b101001111;assign rom[10283] = 'b000111010;assign rom[10284] = 'b101110110;assign rom[10285] = 'b101100010;assign rom[10286] = 'b101001100;assign rom[10287] = 'b001001010;assign rom[10288] = 'b111011010;assign rom[10289] = 'b111011010;assign rom[10290] = 'b111011010;assign rom[10291] = 'b111011010;assign rom[10292] = 'b111011000;assign rom[10293] = 'b111011000;assign rom[10294] = 'b111011000;assign rom[10295] = 'b111011000;assign rom[10296] = 'b101111000;assign rom[10297] = 'b000110011;assign rom[10298] = 'b110000010;assign rom[10299] = 'b001101010;assign rom[10300] = 'b001011000;assign rom[10301] = 'b101001000;assign rom[10302] = 'b000101011;assign rom[10303] = 'b110000010;assign rom[10304] = 'b111000000;assign rom[10305] = 'b101001100;assign rom[10306] = 'b001001010;assign rom[10307] = 'b111111000;assign rom[10308] = 'b111101000;assign rom[10309] = 'b101001111;assign rom[10310] = 'b000111010;assign rom[10311] = 'b101110110;assign rom[10312] = 'b101100010;assign rom[10313] = 'b101001100;assign rom[10314] = 'b001001010;assign rom[10315] = 'b111011010;assign rom[10316] = 'b111011010;assign rom[10317] = 'b111011010;assign rom[10318] = 'b111011010;assign rom[10319] = 'b111011000;assign rom[10320] = 'b111011000;assign rom[10321] = 'b111011000;assign rom[10322] = 'b111011000;assign rom[10323] = 'b101111000;assign rom[10324] = 'b000110011;assign rom[10325] = 'b110000010;assign rom[10326] = 'b001101010;assign rom[10327] = 'b001011000;assign rom[10328] = 'b101001000;assign rom[10329] = 'b000101011;assign rom[10330] = 'b110000010;assign rom[10331] = 'b111000000;assign rom[10332] = 'b101001100;assign rom[10333] = 'b001001010;assign rom[10334] = 'b111111000;assign rom[10335] = 'b111101000;assign rom[10336] = 'b101001111;assign rom[10337] = 'b000111010;assign rom[10338] = 'b101110110;assign rom[10339] = 'b101100010;assign rom[10340] = 'b101001100;assign rom[10341] = 'b001001010;assign rom[10342] = 'b111011010;assign rom[10343] = 'b111011010;assign rom[10344] = 'b111011010;assign rom[10345] = 'b111011010;assign rom[10346] = 'b111011000;assign rom[10347] = 'b111011000;assign rom[10348] = 'b111011000;assign rom[10349] = 'b111011000;assign rom[10350] = 'b101111000;assign rom[10351] = 'b000110011;assign rom[10352] = 'b110000010;assign rom[10353] = 'b001101010;assign rom[10354] = 'b001011000;assign rom[10355] = 'b101001000;assign rom[10356] = 'b000101011;assign rom[10357] = 'b110000010;assign rom[10358] = 'b111000000;assign rom[10359] = 'b101001100;assign rom[10360] = 'b001001010;assign rom[10361] = 'b001000110;assign rom[10362] = 'b001100100;assign rom[10363] = 'b101100010;assign rom[10364] = 'b101001100;assign rom[10365] = 'b001001010;assign rom[10366] = 'b111011010;assign rom[10367] = 'b111011010;assign rom[10368] = 'b111011010;assign rom[10369] = 'b111011010;assign rom[10370] = 'b111011000;assign rom[10371] = 'b111011000;assign rom[10372] = 'b111011000;assign rom[10373] = 'b111011000;assign rom[10374] = 'b101111000;assign rom[10375] = 'b000110011;assign rom[10376] = 'b110000010;assign rom[10377] = 'b001101010;assign rom[10378] = 'b001011000;assign rom[10379] = 'b101001000;assign rom[10380] = 'b000101011;assign rom[10381] = 'b110000010;assign rom[10382] = 'b111000000;assign rom[10383] = 'b101001100;assign rom[10384] = 'b001001010;assign rom[10385] = 'b111111000;assign rom[10386] = 'b111101000;assign rom[10387] = 'b101001111;assign rom[10388] = 'b000111010;assign rom[10389] = 'b101110110;assign rom[10390] = 'b101100010;assign rom[10391] = 'b101001100;assign rom[10392] = 'b001001010;assign rom[10393] = 'b111011010;assign rom[10394] = 'b111011010;assign rom[10395] = 'b111011010;assign rom[10396] = 'b111011010;assign rom[10397] = 'b111011000;assign rom[10398] = 'b111011000;assign rom[10399] = 'b111011000;assign rom[10400] = 'b111011000;assign rom[10401] = 'b101111000;assign rom[10402] = 'b000110011;assign rom[10403] = 'b110000010;assign rom[10404] = 'b001101010;assign rom[10405] = 'b001011000;assign rom[10406] = 'b101001000;assign rom[10407] = 'b000101011;assign rom[10408] = 'b110000010;assign rom[10409] = 'b111000000;assign rom[10410] = 'b101001100;assign rom[10411] = 'b001001010;assign rom[10412] = 'b111111000;assign rom[10413] = 'b111101000;assign rom[10414] = 'b101001111;assign rom[10415] = 'b000111010;assign rom[10416] = 'b101110110;assign rom[10417] = 'b101100010;assign rom[10418] = 'b101001100;assign rom[10419] = 'b001001010;assign rom[10420] = 'b111011010;assign rom[10421] = 'b111011010;assign rom[10422] = 'b111011010;assign rom[10423] = 'b111011010;assign rom[10424] = 'b111011000;assign rom[10425] = 'b111011000;assign rom[10426] = 'b111011000;assign rom[10427] = 'b111011000;assign rom[10428] = 'b101111000;assign rom[10429] = 'b000110011;assign rom[10430] = 'b110000010;assign rom[10431] = 'b001101010;assign rom[10432] = 'b001011000;assign rom[10433] = 'b101001000;assign rom[10434] = 'b000101011;assign rom[10435] = 'b110000010;assign rom[10436] = 'b111000000;assign rom[10437] = 'b101001100;assign rom[10438] = 'b001001010;assign rom[10439] = 'b111111000;assign rom[10440] = 'b111101000;assign rom[10441] = 'b101001111;assign rom[10442] = 'b000111010;assign rom[10443] = 'b101110110;assign rom[10444] = 'b101100010;assign rom[10445] = 'b101001100;assign rom[10446] = 'b001001010;assign rom[10447] = 'b111011010;assign rom[10448] = 'b111011010;assign rom[10449] = 'b111011010;assign rom[10450] = 'b111011010;assign rom[10451] = 'b111011000;assign rom[10452] = 'b111011000;assign rom[10453] = 'b111011000;assign rom[10454] = 'b111011000;assign rom[10455] = 'b101111000;assign rom[10456] = 'b000110011;assign rom[10457] = 'b110000010;assign rom[10458] = 'b001101010;assign rom[10459] = 'b001011000;assign rom[10460] = 'b101001000;assign rom[10461] = 'b000101011;assign rom[10462] = 'b110000010;assign rom[10463] = 'b111000000;assign rom[10464] = 'b101001100;assign rom[10465] = 'b001001010;assign rom[10466] = 'b111111000;assign rom[10467] = 'b111101000;assign rom[10468] = 'b101001111;assign rom[10469] = 'b000111010;assign rom[10470] = 'b101110110;assign rom[10471] = 'b101100010;assign rom[10472] = 'b101001100;assign rom[10473] = 'b001001010;assign rom[10474] = 'b111011010;assign rom[10475] = 'b111011010;assign rom[10476] = 'b111011010;assign rom[10477] = 'b111011010;assign rom[10478] = 'b111011000;assign rom[10479] = 'b111011000;assign rom[10480] = 'b111011000;assign rom[10481] = 'b111011000;assign rom[10482] = 'b101111000;assign rom[10483] = 'b000110011;assign rom[10484] = 'b110000010;assign rom[10485] = 'b001101010;assign rom[10486] = 'b001011000;assign rom[10487] = 'b101001000;assign rom[10488] = 'b000101011;assign rom[10489] = 'b110000010;assign rom[10490] = 'b111000000;assign rom[10491] = 'b101001100;assign rom[10492] = 'b001001010;assign rom[10493] = 'b111111000;assign rom[10494] = 'b111101000;assign rom[10495] = 'b101001111;assign rom[10496] = 'b000111010;assign rom[10497] = 'b101110110;assign rom[10498] = 'b101100010;assign rom[10499] = 'b101001100;assign rom[10500] = 'b001001010;assign rom[10501] = 'b111011010;assign rom[10502] = 'b111011010;assign rom[10503] = 'b111011010;assign rom[10504] = 'b111011010;assign rom[10505] = 'b111011000;assign rom[10506] = 'b111011000;assign rom[10507] = 'b111011000;assign rom[10508] = 'b111011000;assign rom[10509] = 'b101111000;assign rom[10510] = 'b000110011;assign rom[10511] = 'b110000010;assign rom[10512] = 'b001101010;assign rom[10513] = 'b001011000;assign rom[10514] = 'b101001000;assign rom[10515] = 'b000101011;assign rom[10516] = 'b110000010;assign rom[10517] = 'b111000000;assign rom[10518] = 'b101001100;assign rom[10519] = 'b001001010;assign rom[10520] = 'b111111000;assign rom[10521] = 'b111101000;assign rom[10522] = 'b101001111;assign rom[10523] = 'b000111010;assign rom[10524] = 'b101110110;assign rom[10525] = 'b101100010;assign rom[10526] = 'b101001100;assign rom[10527] = 'b001001010;assign rom[10528] = 'b111011010;assign rom[10529] = 'b111011010;assign rom[10530] = 'b111011010;assign rom[10531] = 'b111011010;assign rom[10532] = 'b111011000;assign rom[10533] = 'b111011000;assign rom[10534] = 'b111011000;assign rom[10535] = 'b111011000;assign rom[10536] = 'b101111000;assign rom[10537] = 'b000110011;assign rom[10538] = 'b110000010;assign rom[10539] = 'b001101010;assign rom[10540] = 'b001011000;assign rom[10541] = 'b101001000;assign rom[10542] = 'b000101011;assign rom[10543] = 'b110000010;assign rom[10544] = 'b111000000;assign rom[10545] = 'b101001100;assign rom[10546] = 'b001001010;assign rom[10547] = 'b111111000;assign rom[10548] = 'b111101000;assign rom[10549] = 'b101001111;assign rom[10550] = 'b000111010;assign rom[10551] = 'b101110110;assign rom[10552] = 'b101100010;assign rom[10553] = 'b101001100;assign rom[10554] = 'b001001010;assign rom[10555] = 'b111011010;assign rom[10556] = 'b111011010;assign rom[10557] = 'b111011010;assign rom[10558] = 'b111011010;assign rom[10559] = 'b111011000;assign rom[10560] = 'b111011000;assign rom[10561] = 'b111011000;assign rom[10562] = 'b111011000;assign rom[10563] = 'b101111000;assign rom[10564] = 'b000110011;assign rom[10565] = 'b110000010;assign rom[10566] = 'b001101010;assign rom[10567] = 'b001011000;assign rom[10568] = 'b101001000;assign rom[10569] = 'b000101011;assign rom[10570] = 'b110000010;assign rom[10571] = 'b111000000;assign rom[10572] = 'b101001100;assign rom[10573] = 'b001001010;assign rom[10574] = 'b111111000;assign rom[10575] = 'b111101000;assign rom[10576] = 'b101001111;assign rom[10577] = 'b000111010;assign rom[10578] = 'b101110110;assign rom[10579] = 'b101100010;assign rom[10580] = 'b101001100;assign rom[10581] = 'b001001010;assign rom[10582] = 'b111011010;assign rom[10583] = 'b111011010;assign rom[10584] = 'b111011010;assign rom[10585] = 'b111011010;assign rom[10586] = 'b111011000;assign rom[10587] = 'b111011000;assign rom[10588] = 'b111011000;assign rom[10589] = 'b111011000;assign rom[10590] = 'b101111000;assign rom[10591] = 'b000110011;assign rom[10592] = 'b110000010;assign rom[10593] = 'b001101010;assign rom[10594] = 'b001011000;assign rom[10595] = 'b101001000;assign rom[10596] = 'b000101011;assign rom[10597] = 'b110000010;assign rom[10598] = 'b111000000;assign rom[10599] = 'b101001100;assign rom[10600] = 'b001001010;assign rom[10601] = 'b001000110;assign rom[10602] = 'b001100100;assign rom[10603] = 'b101100010;assign rom[10604] = 'b101001100;assign rom[10605] = 'b001001010;assign rom[10606] = 'b111011010;assign rom[10607] = 'b111011010;assign rom[10608] = 'b111011010;assign rom[10609] = 'b111011010;assign rom[10610] = 'b111011000;assign rom[10611] = 'b111011000;assign rom[10612] = 'b111011000;assign rom[10613] = 'b111011000;assign rom[10614] = 'b101111000;assign rom[10615] = 'b000110011;assign rom[10616] = 'b110000010;assign rom[10617] = 'b001101010;assign rom[10618] = 'b001011000;assign rom[10619] = 'b101001000;assign rom[10620] = 'b000101011;assign rom[10621] = 'b110000010;assign rom[10622] = 'b111000000;assign rom[10623] = 'b101001100;assign rom[10624] = 'b001001010;assign rom[10625] = 'b111111000;assign rom[10626] = 'b111101000;assign rom[10627] = 'b101001111;assign rom[10628] = 'b000111010;assign rom[10629] = 'b101110110;assign rom[10630] = 'b101100010;assign rom[10631] = 'b101001100;assign rom[10632] = 'b001001010;assign rom[10633] = 'b111011010;assign rom[10634] = 'b111011010;assign rom[10635] = 'b111011010;assign rom[10636] = 'b111011010;assign rom[10637] = 'b111011000;assign rom[10638] = 'b111011000;assign rom[10639] = 'b111011000;assign rom[10640] = 'b111011000;assign rom[10641] = 'b101111000;assign rom[10642] = 'b000110011;assign rom[10643] = 'b110000010;assign rom[10644] = 'b001101010;assign rom[10645] = 'b001011000;assign rom[10646] = 'b101001000;assign rom[10647] = 'b000101011;assign rom[10648] = 'b110000010;assign rom[10649] = 'b111000000;assign rom[10650] = 'b101001100;assign rom[10651] = 'b001001010;assign rom[10652] = 'b111111000;assign rom[10653] = 'b111101000;assign rom[10654] = 'b101001111;assign rom[10655] = 'b000111010;assign rom[10656] = 'b101110110;assign rom[10657] = 'b101100010;assign rom[10658] = 'b101001100;assign rom[10659] = 'b001001010;assign rom[10660] = 'b111011010;assign rom[10661] = 'b111011010;assign rom[10662] = 'b111011010;assign rom[10663] = 'b111011010;assign rom[10664] = 'b111011000;assign rom[10665] = 'b111011000;assign rom[10666] = 'b111011000;assign rom[10667] = 'b111011000;assign rom[10668] = 'b101111000;assign rom[10669] = 'b000110011;assign rom[10670] = 'b110000010;assign rom[10671] = 'b001101010;assign rom[10672] = 'b001011000;assign rom[10673] = 'b101001000;assign rom[10674] = 'b000101011;assign rom[10675] = 'b110000010;assign rom[10676] = 'b111000000;assign rom[10677] = 'b101001100;assign rom[10678] = 'b001001010;assign rom[10679] = 'b111111000;assign rom[10680] = 'b111101000;assign rom[10681] = 'b101001111;assign rom[10682] = 'b000111010;assign rom[10683] = 'b101110110;assign rom[10684] = 'b101100010;assign rom[10685] = 'b101001100;assign rom[10686] = 'b001001010;assign rom[10687] = 'b111011010;assign rom[10688] = 'b111011010;assign rom[10689] = 'b111011010;assign rom[10690] = 'b111011010;assign rom[10691] = 'b111011000;assign rom[10692] = 'b111011000;assign rom[10693] = 'b111011000;assign rom[10694] = 'b111011000;assign rom[10695] = 'b101111000;assign rom[10696] = 'b000110011;assign rom[10697] = 'b110000010;assign rom[10698] = 'b001101010;assign rom[10699] = 'b001011000;assign rom[10700] = 'b101001000;assign rom[10701] = 'b000101011;assign rom[10702] = 'b110000010;assign rom[10703] = 'b111000000;assign rom[10704] = 'b101001100;assign rom[10705] = 'b001001010;assign rom[10706] = 'b111111000;assign rom[10707] = 'b111101000;assign rom[10708] = 'b101001111;assign rom[10709] = 'b000111010;assign rom[10710] = 'b101110110;assign rom[10711] = 'b101100010;assign rom[10712] = 'b101001100;assign rom[10713] = 'b001001010;assign rom[10714] = 'b111011010;assign rom[10715] = 'b111011010;assign rom[10716] = 'b111011010;assign rom[10717] = 'b111011010;assign rom[10718] = 'b111011000;assign rom[10719] = 'b111011000;assign rom[10720] = 'b111011000;assign rom[10721] = 'b111011000;assign rom[10722] = 'b101111000;assign rom[10723] = 'b000110011;assign rom[10724] = 'b110000010;assign rom[10725] = 'b001101010;assign rom[10726] = 'b001011000;assign rom[10727] = 'b101001000;assign rom[10728] = 'b000101011;assign rom[10729] = 'b110000010;assign rom[10730] = 'b111000000;assign rom[10731] = 'b101001100;assign rom[10732] = 'b001001010;assign rom[10733] = 'b111111000;assign rom[10734] = 'b111101000;assign rom[10735] = 'b101001111;assign rom[10736] = 'b000111010;assign rom[10737] = 'b101110110;assign rom[10738] = 'b101100010;assign rom[10739] = 'b101001100;assign rom[10740] = 'b001001010;assign rom[10741] = 'b111011010;assign rom[10742] = 'b111011010;assign rom[10743] = 'b111011010;assign rom[10744] = 'b111011010;assign rom[10745] = 'b111011000;assign rom[10746] = 'b111011000;assign rom[10747] = 'b111011000;assign rom[10748] = 'b111011000;assign rom[10749] = 'b101111000;assign rom[10750] = 'b000110011;assign rom[10751] = 'b110000010;assign rom[10752] = 'b001101010;assign rom[10753] = 'b001011000;assign rom[10754] = 'b101001000;assign rom[10755] = 'b000101011;assign rom[10756] = 'b110000010;assign rom[10757] = 'b111000000;assign rom[10758] = 'b101001100;assign rom[10759] = 'b001001010;assign rom[10760] = 'b111111000;assign rom[10761] = 'b111101000;assign rom[10762] = 'b101001111;assign rom[10763] = 'b000111010;assign rom[10764] = 'b101110110;assign rom[10765] = 'b101100010;assign rom[10766] = 'b101001100;assign rom[10767] = 'b001001010;assign rom[10768] = 'b111011010;assign rom[10769] = 'b111011010;assign rom[10770] = 'b111011010;assign rom[10771] = 'b111011010;assign rom[10772] = 'b111011000;assign rom[10773] = 'b111011000;assign rom[10774] = 'b111011000;assign rom[10775] = 'b111011000;assign rom[10776] = 'b101111000;assign rom[10777] = 'b000110011;assign rom[10778] = 'b110000010;assign rom[10779] = 'b001101010;assign rom[10780] = 'b001011000;assign rom[10781] = 'b101001000;assign rom[10782] = 'b000101011;assign rom[10783] = 'b110000010;assign rom[10784] = 'b111000000;assign rom[10785] = 'b101001100;assign rom[10786] = 'b001001010;assign rom[10787] = 'b111111000;assign rom[10788] = 'b111101000;assign rom[10789] = 'b101001111;assign rom[10790] = 'b000111010;assign rom[10791] = 'b101110110;assign rom[10792] = 'b101100010;assign rom[10793] = 'b101001100;assign rom[10794] = 'b001001010;assign rom[10795] = 'b111011010;assign rom[10796] = 'b111011010;assign rom[10797] = 'b111011010;assign rom[10798] = 'b111011010;assign rom[10799] = 'b111011000;assign rom[10800] = 'b111011000;assign rom[10801] = 'b111011000;assign rom[10802] = 'b111011000;assign rom[10803] = 'b101111000;assign rom[10804] = 'b000110011;assign rom[10805] = 'b110000010;assign rom[10806] = 'b001101010;assign rom[10807] = 'b001011000;assign rom[10808] = 'b101001000;assign rom[10809] = 'b000101011;assign rom[10810] = 'b110000010;assign rom[10811] = 'b111000000;assign rom[10812] = 'b101001100;assign rom[10813] = 'b001001010;assign rom[10814] = 'b111111000;assign rom[10815] = 'b111101000;assign rom[10816] = 'b101001111;assign rom[10817] = 'b000111010;assign rom[10818] = 'b101110110;assign rom[10819] = 'b101100010;assign rom[10820] = 'b101001100;assign rom[10821] = 'b001001010;assign rom[10822] = 'b111011010;assign rom[10823] = 'b111011010;assign rom[10824] = 'b111011010;assign rom[10825] = 'b111011010;assign rom[10826] = 'b111011000;assign rom[10827] = 'b111011000;assign rom[10828] = 'b111011000;assign rom[10829] = 'b111011000;assign rom[10830] = 'b101111000;assign rom[10831] = 'b000110011;assign rom[10832] = 'b110000010;assign rom[10833] = 'b001101010;assign rom[10834] = 'b001011000;assign rom[10835] = 'b101001000;assign rom[10836] = 'b000101011;assign rom[10837] = 'b110000010;assign rom[10838] = 'b111000000;assign rom[10839] = 'b101001100;assign rom[10840] = 'b001001010;assign rom[10841] = 'b001000110;assign rom[10842] = 'b001100100;assign rom[10843] = 'b101100010;assign rom[10844] = 'b101001100;assign rom[10845] = 'b001001010;assign rom[10846] = 'b111011010;assign rom[10847] = 'b111011010;assign rom[10848] = 'b111011010;assign rom[10849] = 'b111011010;assign rom[10850] = 'b111011000;assign rom[10851] = 'b111011000;assign rom[10852] = 'b111011000;assign rom[10853] = 'b111011000;assign rom[10854] = 'b101111000;assign rom[10855] = 'b000110011;assign rom[10856] = 'b110000010;assign rom[10857] = 'b001101010;assign rom[10858] = 'b001011000;assign rom[10859] = 'b101001000;assign rom[10860] = 'b000101011;assign rom[10861] = 'b110000010;assign rom[10862] = 'b111000000;assign rom[10863] = 'b101001100;assign rom[10864] = 'b001001010;assign rom[10865] = 'b111111000;assign rom[10866] = 'b111101000;assign rom[10867] = 'b101001111;assign rom[10868] = 'b000111010;assign rom[10869] = 'b101110110;assign rom[10870] = 'b101100010;assign rom[10871] = 'b101001100;assign rom[10872] = 'b001001010;assign rom[10873] = 'b111011010;assign rom[10874] = 'b111011010;assign rom[10875] = 'b111011010;assign rom[10876] = 'b111011010;assign rom[10877] = 'b111011000;assign rom[10878] = 'b111011000;assign rom[10879] = 'b111011000;assign rom[10880] = 'b111011000;assign rom[10881] = 'b101111000;assign rom[10882] = 'b000110011;assign rom[10883] = 'b110000010;assign rom[10884] = 'b001101010;assign rom[10885] = 'b001011000;assign rom[10886] = 'b101001000;assign rom[10887] = 'b000101011;assign rom[10888] = 'b110000010;assign rom[10889] = 'b111000000;assign rom[10890] = 'b101001100;assign rom[10891] = 'b001001010;assign rom[10892] = 'b111111000;assign rom[10893] = 'b111101000;assign rom[10894] = 'b101001111;assign rom[10895] = 'b000111010;assign rom[10896] = 'b101110110;assign rom[10897] = 'b101100010;assign rom[10898] = 'b101001100;assign rom[10899] = 'b001001010;assign rom[10900] = 'b111011010;assign rom[10901] = 'b111011010;assign rom[10902] = 'b111011010;assign rom[10903] = 'b111011010;assign rom[10904] = 'b111011000;assign rom[10905] = 'b111011000;assign rom[10906] = 'b111011000;assign rom[10907] = 'b111011000;assign rom[10908] = 'b101111000;assign rom[10909] = 'b000110011;assign rom[10910] = 'b110000010;assign rom[10911] = 'b001101010;assign rom[10912] = 'b001011000;assign rom[10913] = 'b101001000;assign rom[10914] = 'b000101011;assign rom[10915] = 'b110000010;assign rom[10916] = 'b111000000;assign rom[10917] = 'b101001100;assign rom[10918] = 'b001001010;assign rom[10919] = 'b111111000;assign rom[10920] = 'b111101000;assign rom[10921] = 'b101001111;assign rom[10922] = 'b000111010;assign rom[10923] = 'b101110110;assign rom[10924] = 'b101100010;assign rom[10925] = 'b101001100;assign rom[10926] = 'b001001010;assign rom[10927] = 'b111011010;assign rom[10928] = 'b111011010;assign rom[10929] = 'b111011010;assign rom[10930] = 'b111011010;assign rom[10931] = 'b111011000;assign rom[10932] = 'b111011000;assign rom[10933] = 'b111011000;assign rom[10934] = 'b111011000;assign rom[10935] = 'b101111000;assign rom[10936] = 'b000110011;assign rom[10937] = 'b110000010;assign rom[10938] = 'b001101010;assign rom[10939] = 'b001011000;assign rom[10940] = 'b101001000;assign rom[10941] = 'b000101011;assign rom[10942] = 'b110000010;assign rom[10943] = 'b111000000;assign rom[10944] = 'b101001100;assign rom[10945] = 'b001001010;assign rom[10946] = 'b111111000;assign rom[10947] = 'b111101000;assign rom[10948] = 'b101001111;assign rom[10949] = 'b000111010;assign rom[10950] = 'b101110110;assign rom[10951] = 'b101100010;assign rom[10952] = 'b101001100;assign rom[10953] = 'b001001010;assign rom[10954] = 'b111011010;assign rom[10955] = 'b111011010;assign rom[10956] = 'b111011010;assign rom[10957] = 'b111011010;assign rom[10958] = 'b111011000;assign rom[10959] = 'b111011000;assign rom[10960] = 'b111011000;assign rom[10961] = 'b111011000;assign rom[10962] = 'b101111000;assign rom[10963] = 'b000110011;assign rom[10964] = 'b110000010;assign rom[10965] = 'b001101010;assign rom[10966] = 'b001011000;assign rom[10967] = 'b101001000;assign rom[10968] = 'b000101011;assign rom[10969] = 'b110000010;assign rom[10970] = 'b111000000;assign rom[10971] = 'b101001100;assign rom[10972] = 'b001001010;assign rom[10973] = 'b111111000;assign rom[10974] = 'b111101000;assign rom[10975] = 'b101001111;assign rom[10976] = 'b000111010;assign rom[10977] = 'b101110110;assign rom[10978] = 'b101100010;assign rom[10979] = 'b101001100;assign rom[10980] = 'b001001010;assign rom[10981] = 'b111011010;assign rom[10982] = 'b111011010;assign rom[10983] = 'b111011010;assign rom[10984] = 'b111011010;assign rom[10985] = 'b111011000;assign rom[10986] = 'b111011000;assign rom[10987] = 'b111011000;assign rom[10988] = 'b111011000;assign rom[10989] = 'b101111000;assign rom[10990] = 'b000110011;assign rom[10991] = 'b110000010;assign rom[10992] = 'b001101010;assign rom[10993] = 'b001011000;assign rom[10994] = 'b101001000;assign rom[10995] = 'b000101011;assign rom[10996] = 'b110000010;assign rom[10997] = 'b111000000;assign rom[10998] = 'b101001100;assign rom[10999] = 'b001001010;assign rom[11000] = 'b111111000;assign rom[11001] = 'b111101000;assign rom[11002] = 'b101001111;assign rom[11003] = 'b000111010;assign rom[11004] = 'b101110110;assign rom[11005] = 'b101100010;assign rom[11006] = 'b101001100;assign rom[11007] = 'b001001010;assign rom[11008] = 'b111011010;assign rom[11009] = 'b111011010;assign rom[11010] = 'b111011010;assign rom[11011] = 'b111011010;assign rom[11012] = 'b111011000;assign rom[11013] = 'b111011000;assign rom[11014] = 'b111011000;assign rom[11015] = 'b111011000;assign rom[11016] = 'b101111000;assign rom[11017] = 'b000110011;assign rom[11018] = 'b110000010;assign rom[11019] = 'b001101010;assign rom[11020] = 'b001011000;assign rom[11021] = 'b101001000;assign rom[11022] = 'b000101011;assign rom[11023] = 'b110000010;assign rom[11024] = 'b111000000;assign rom[11025] = 'b101001100;assign rom[11026] = 'b001001010;assign rom[11027] = 'b111111000;assign rom[11028] = 'b111101000;assign rom[11029] = 'b101001111;assign rom[11030] = 'b000111010;assign rom[11031] = 'b101110110;assign rom[11032] = 'b101100010;assign rom[11033] = 'b101001100;assign rom[11034] = 'b001001010;assign rom[11035] = 'b111011010;assign rom[11036] = 'b111011010;assign rom[11037] = 'b111011010;assign rom[11038] = 'b111011010;assign rom[11039] = 'b111011000;assign rom[11040] = 'b111011000;assign rom[11041] = 'b111011000;assign rom[11042] = 'b111011000;assign rom[11043] = 'b101111000;assign rom[11044] = 'b000110011;assign rom[11045] = 'b110000010;assign rom[11046] = 'b001101010;assign rom[11047] = 'b001011000;assign rom[11048] = 'b101001000;assign rom[11049] = 'b000101011;assign rom[11050] = 'b110000010;assign rom[11051] = 'b111000000;assign rom[11052] = 'b101001100;assign rom[11053] = 'b001001010;assign rom[11054] = 'b111111000;assign rom[11055] = 'b111101000;assign rom[11056] = 'b101001111;assign rom[11057] = 'b000111010;assign rom[11058] = 'b101110110;assign rom[11059] = 'b101100010;assign rom[11060] = 'b101001100;assign rom[11061] = 'b001001010;assign rom[11062] = 'b111011010;assign rom[11063] = 'b111011010;assign rom[11064] = 'b111011010;assign rom[11065] = 'b111011010;assign rom[11066] = 'b111011000;assign rom[11067] = 'b111011000;assign rom[11068] = 'b111011000;assign rom[11069] = 'b111011000;assign rom[11070] = 'b101111000;assign rom[11071] = 'b000110011;assign rom[11072] = 'b110000010;assign rom[11073] = 'b001101010;assign rom[11074] = 'b001011000;assign rom[11075] = 'b101001000;assign rom[11076] = 'b000101011;assign rom[11077] = 'b110000010;assign rom[11078] = 'b111000000;assign rom[11079] = 'b101001100;assign rom[11080] = 'b001001010;assign rom[11081] = 'b001000110;assign rom[11082] = 'b001100100;assign rom[11083] = 'b101100010;assign rom[11084] = 'b101001100;assign rom[11085] = 'b001001010;assign rom[11086] = 'b111011010;assign rom[11087] = 'b111011010;assign rom[11088] = 'b111011010;assign rom[11089] = 'b111011010;assign rom[11090] = 'b111011000;assign rom[11091] = 'b111011000;assign rom[11092] = 'b111011000;assign rom[11093] = 'b111011000;assign rom[11094] = 'b101111000;assign rom[11095] = 'b000110011;assign rom[11096] = 'b110000010;assign rom[11097] = 'b001101010;assign rom[11098] = 'b001011000;assign rom[11099] = 'b101001000;assign rom[11100] = 'b000101011;assign rom[11101] = 'b110000010;assign rom[11102] = 'b111000000;assign rom[11103] = 'b101001100;assign rom[11104] = 'b001001010;assign rom[11105] = 'b111111000;assign rom[11106] = 'b111101000;assign rom[11107] = 'b101001111;assign rom[11108] = 'b000111010;assign rom[11109] = 'b101110110;assign rom[11110] = 'b101100010;assign rom[11111] = 'b101001100;assign rom[11112] = 'b001001010;assign rom[11113] = 'b111011010;assign rom[11114] = 'b111011010;assign rom[11115] = 'b111011010;assign rom[11116] = 'b111011010;assign rom[11117] = 'b111011000;assign rom[11118] = 'b111011000;assign rom[11119] = 'b111011000;assign rom[11120] = 'b111011000;assign rom[11121] = 'b101111000;assign rom[11122] = 'b000110011;assign rom[11123] = 'b110000010;assign rom[11124] = 'b001101010;assign rom[11125] = 'b001011000;assign rom[11126] = 'b101001000;assign rom[11127] = 'b000101011;assign rom[11128] = 'b110000010;assign rom[11129] = 'b111000000;assign rom[11130] = 'b101001100;assign rom[11131] = 'b001001010;assign rom[11132] = 'b111111000;assign rom[11133] = 'b111101000;assign rom[11134] = 'b101001111;assign rom[11135] = 'b000111010;assign rom[11136] = 'b101110110;assign rom[11137] = 'b101100010;assign rom[11138] = 'b101001100;assign rom[11139] = 'b001001010;assign rom[11140] = 'b111011010;assign rom[11141] = 'b111011010;assign rom[11142] = 'b111011010;assign rom[11143] = 'b111011010;assign rom[11144] = 'b111011000;assign rom[11145] = 'b111011000;assign rom[11146] = 'b111011000;assign rom[11147] = 'b111011000;assign rom[11148] = 'b101111000;assign rom[11149] = 'b000110011;assign rom[11150] = 'b110000010;assign rom[11151] = 'b001101010;assign rom[11152] = 'b001011000;assign rom[11153] = 'b101001000;assign rom[11154] = 'b000101011;assign rom[11155] = 'b110000010;assign rom[11156] = 'b111000000;assign rom[11157] = 'b101001100;assign rom[11158] = 'b001001010;assign rom[11159] = 'b111111000;assign rom[11160] = 'b111101000;assign rom[11161] = 'b101001111;assign rom[11162] = 'b000111010;assign rom[11163] = 'b101110110;assign rom[11164] = 'b101100010;assign rom[11165] = 'b101001100;assign rom[11166] = 'b001001010;assign rom[11167] = 'b111011010;assign rom[11168] = 'b111011010;assign rom[11169] = 'b111011010;assign rom[11170] = 'b111011010;assign rom[11171] = 'b111011000;assign rom[11172] = 'b111011000;assign rom[11173] = 'b111011000;assign rom[11174] = 'b111011000;assign rom[11175] = 'b101111000;assign rom[11176] = 'b000110011;assign rom[11177] = 'b110000010;assign rom[11178] = 'b001101010;assign rom[11179] = 'b001011000;assign rom[11180] = 'b101001000;assign rom[11181] = 'b000101011;assign rom[11182] = 'b110000010;assign rom[11183] = 'b111000000;assign rom[11184] = 'b101001100;assign rom[11185] = 'b001001010;assign rom[11186] = 'b111111000;assign rom[11187] = 'b111101000;assign rom[11188] = 'b101001111;assign rom[11189] = 'b000111010;assign rom[11190] = 'b101110110;assign rom[11191] = 'b101100010;assign rom[11192] = 'b101001100;assign rom[11193] = 'b001001010;assign rom[11194] = 'b111011010;assign rom[11195] = 'b111011010;assign rom[11196] = 'b111011010;assign rom[11197] = 'b111011010;assign rom[11198] = 'b111011000;assign rom[11199] = 'b111011000;assign rom[11200] = 'b111011000;assign rom[11201] = 'b111011000;assign rom[11202] = 'b101111000;assign rom[11203] = 'b000110011;assign rom[11204] = 'b110000010;assign rom[11205] = 'b001101010;assign rom[11206] = 'b001011000;assign rom[11207] = 'b101001000;assign rom[11208] = 'b000101011;assign rom[11209] = 'b110000010;assign rom[11210] = 'b111000000;assign rom[11211] = 'b101001100;assign rom[11212] = 'b001001010;assign rom[11213] = 'b111111000;assign rom[11214] = 'b111101000;assign rom[11215] = 'b101001111;assign rom[11216] = 'b000111010;assign rom[11217] = 'b101110110;assign rom[11218] = 'b101100010;assign rom[11219] = 'b101001100;assign rom[11220] = 'b001001010;assign rom[11221] = 'b111011010;assign rom[11222] = 'b111011010;assign rom[11223] = 'b111011010;assign rom[11224] = 'b111011010;assign rom[11225] = 'b111011000;assign rom[11226] = 'b111011000;assign rom[11227] = 'b111011000;assign rom[11228] = 'b111011000;assign rom[11229] = 'b101111000;assign rom[11230] = 'b000110011;assign rom[11231] = 'b110000010;assign rom[11232] = 'b001101010;assign rom[11233] = 'b001011000;assign rom[11234] = 'b101001000;assign rom[11235] = 'b000101011;assign rom[11236] = 'b110000010;assign rom[11237] = 'b111000000;assign rom[11238] = 'b101001100;assign rom[11239] = 'b001001010;assign rom[11240] = 'b111111000;assign rom[11241] = 'b111101000;assign rom[11242] = 'b101001111;assign rom[11243] = 'b000111010;assign rom[11244] = 'b101110110;assign rom[11245] = 'b101100010;assign rom[11246] = 'b101001100;assign rom[11247] = 'b001001010;assign rom[11248] = 'b111011010;assign rom[11249] = 'b111011010;assign rom[11250] = 'b111011010;assign rom[11251] = 'b111011010;assign rom[11252] = 'b111011000;assign rom[11253] = 'b111011000;assign rom[11254] = 'b111011000;assign rom[11255] = 'b111011000;assign rom[11256] = 'b101111000;assign rom[11257] = 'b000110011;assign rom[11258] = 'b110000010;assign rom[11259] = 'b001101010;assign rom[11260] = 'b001011000;assign rom[11261] = 'b101001000;assign rom[11262] = 'b000101011;assign rom[11263] = 'b110000010;assign rom[11264] = 'b111000000;assign rom[11265] = 'b101001100;assign rom[11266] = 'b001001010;assign rom[11267] = 'b111111000;assign rom[11268] = 'b111101000;assign rom[11269] = 'b101001111;assign rom[11270] = 'b000111010;assign rom[11271] = 'b101110110;assign rom[11272] = 'b101100010;assign rom[11273] = 'b101001100;assign rom[11274] = 'b001001010;assign rom[11275] = 'b111011010;assign rom[11276] = 'b111011010;assign rom[11277] = 'b111011010;assign rom[11278] = 'b111011010;assign rom[11279] = 'b111011000;assign rom[11280] = 'b111011000;assign rom[11281] = 'b111011000;assign rom[11282] = 'b111011000;assign rom[11283] = 'b101111000;assign rom[11284] = 'b000110011;assign rom[11285] = 'b110000010;assign rom[11286] = 'b001101010;assign rom[11287] = 'b001011000;assign rom[11288] = 'b101001000;assign rom[11289] = 'b000101011;assign rom[11290] = 'b110000010;assign rom[11291] = 'b111000000;assign rom[11292] = 'b101001100;assign rom[11293] = 'b001001010;assign rom[11294] = 'b111111000;assign rom[11295] = 'b111101000;assign rom[11296] = 'b101001111;assign rom[11297] = 'b000111010;assign rom[11298] = 'b101110110;assign rom[11299] = 'b101100010;assign rom[11300] = 'b101001100;assign rom[11301] = 'b001001010;assign rom[11302] = 'b111011010;assign rom[11303] = 'b111011010;assign rom[11304] = 'b111011010;assign rom[11305] = 'b111011010;assign rom[11306] = 'b111011000;assign rom[11307] = 'b111011000;assign rom[11308] = 'b111011000;assign rom[11309] = 'b111011000;assign rom[11310] = 'b101111000;assign rom[11311] = 'b000110011;assign rom[11312] = 'b110000010;assign rom[11313] = 'b001101010;assign rom[11314] = 'b001011000;assign rom[11315] = 'b101001000;assign rom[11316] = 'b000101011;assign rom[11317] = 'b110000010;assign rom[11318] = 'b111000000;assign rom[11319] = 'b101001100;assign rom[11320] = 'b001001010;assign rom[11321] = 'b001000110;assign rom[11322] = 'b001100100;assign rom[11323] = 'b101100010;assign rom[11324] = 'b101001100;assign rom[11325] = 'b001001010;assign rom[11326] = 'b111011010;assign rom[11327] = 'b111011010;assign rom[11328] = 'b111011010;assign rom[11329] = 'b111011010;assign rom[11330] = 'b111011000;assign rom[11331] = 'b111011000;assign rom[11332] = 'b111011000;assign rom[11333] = 'b111011000;assign rom[11334] = 'b101111000;assign rom[11335] = 'b000110011;assign rom[11336] = 'b110000010;assign rom[11337] = 'b001101010;assign rom[11338] = 'b001011000;assign rom[11339] = 'b101001000;assign rom[11340] = 'b000101011;assign rom[11341] = 'b110000010;assign rom[11342] = 'b111000000;assign rom[11343] = 'b101001100;assign rom[11344] = 'b001001010;assign rom[11345] = 'b111111000;assign rom[11346] = 'b111101000;assign rom[11347] = 'b101001111;assign rom[11348] = 'b000111010;assign rom[11349] = 'b101110110;assign rom[11350] = 'b101100010;assign rom[11351] = 'b101001100;assign rom[11352] = 'b001001010;assign rom[11353] = 'b111011010;assign rom[11354] = 'b111011010;assign rom[11355] = 'b111011010;assign rom[11356] = 'b111011010;assign rom[11357] = 'b111011000;assign rom[11358] = 'b111011000;assign rom[11359] = 'b111011000;assign rom[11360] = 'b111011000;assign rom[11361] = 'b101111000;assign rom[11362] = 'b000110011;assign rom[11363] = 'b110000010;assign rom[11364] = 'b001101010;assign rom[11365] = 'b001011000;assign rom[11366] = 'b101001000;assign rom[11367] = 'b000101011;assign rom[11368] = 'b110000010;assign rom[11369] = 'b111000000;assign rom[11370] = 'b101001100;assign rom[11371] = 'b001001010;assign rom[11372] = 'b111111000;assign rom[11373] = 'b111101000;assign rom[11374] = 'b101001111;assign rom[11375] = 'b000111010;assign rom[11376] = 'b101110110;assign rom[11377] = 'b101100010;assign rom[11378] = 'b101001100;assign rom[11379] = 'b001001010;assign rom[11380] = 'b111011010;assign rom[11381] = 'b111011010;assign rom[11382] = 'b111011010;assign rom[11383] = 'b111011010;assign rom[11384] = 'b111011000;assign rom[11385] = 'b111011000;assign rom[11386] = 'b111011000;assign rom[11387] = 'b111011000;assign rom[11388] = 'b101111000;assign rom[11389] = 'b000110011;assign rom[11390] = 'b110000010;assign rom[11391] = 'b001101010;assign rom[11392] = 'b001011000;assign rom[11393] = 'b101001000;assign rom[11394] = 'b000101011;assign rom[11395] = 'b110000010;assign rom[11396] = 'b111000000;assign rom[11397] = 'b101001100;assign rom[11398] = 'b001001010;assign rom[11399] = 'b111111000;assign rom[11400] = 'b111101000;assign rom[11401] = 'b101001111;assign rom[11402] = 'b000111010;assign rom[11403] = 'b101110110;assign rom[11404] = 'b101100010;assign rom[11405] = 'b101001100;assign rom[11406] = 'b001001010;assign rom[11407] = 'b111011010;assign rom[11408] = 'b111011010;assign rom[11409] = 'b111011010;assign rom[11410] = 'b111011010;assign rom[11411] = 'b111011000;assign rom[11412] = 'b111011000;assign rom[11413] = 'b111011000;assign rom[11414] = 'b111011000;assign rom[11415] = 'b101111000;assign rom[11416] = 'b000110011;assign rom[11417] = 'b110000010;assign rom[11418] = 'b001101010;assign rom[11419] = 'b001011000;assign rom[11420] = 'b101001000;assign rom[11421] = 'b000101011;assign rom[11422] = 'b110000010;assign rom[11423] = 'b111000000;assign rom[11424] = 'b101001100;assign rom[11425] = 'b001001010;assign rom[11426] = 'b111111000;assign rom[11427] = 'b111101000;assign rom[11428] = 'b101001111;assign rom[11429] = 'b000111010;assign rom[11430] = 'b101110110;assign rom[11431] = 'b101100010;assign rom[11432] = 'b101001100;assign rom[11433] = 'b001001010;assign rom[11434] = 'b111011010;assign rom[11435] = 'b111011010;assign rom[11436] = 'b111011010;assign rom[11437] = 'b111011010;assign rom[11438] = 'b111011000;assign rom[11439] = 'b111011000;assign rom[11440] = 'b111011000;assign rom[11441] = 'b111011000;assign rom[11442] = 'b101111000;assign rom[11443] = 'b000110011;assign rom[11444] = 'b110000010;assign rom[11445] = 'b001101010;assign rom[11446] = 'b001011000;assign rom[11447] = 'b101001000;assign rom[11448] = 'b000101011;assign rom[11449] = 'b110000010;assign rom[11450] = 'b111000000;assign rom[11451] = 'b101001100;assign rom[11452] = 'b001001010;assign rom[11453] = 'b111111000;assign rom[11454] = 'b111101000;assign rom[11455] = 'b101001111;assign rom[11456] = 'b000111010;assign rom[11457] = 'b101110110;assign rom[11458] = 'b101100010;assign rom[11459] = 'b101001100;assign rom[11460] = 'b001001010;assign rom[11461] = 'b111011010;assign rom[11462] = 'b111011010;assign rom[11463] = 'b111011010;assign rom[11464] = 'b111011010;assign rom[11465] = 'b111011000;assign rom[11466] = 'b111011000;assign rom[11467] = 'b111011000;assign rom[11468] = 'b111011000;assign rom[11469] = 'b101111000;assign rom[11470] = 'b000110011;assign rom[11471] = 'b110000010;assign rom[11472] = 'b001101010;assign rom[11473] = 'b001011000;assign rom[11474] = 'b101001000;assign rom[11475] = 'b000101011;assign rom[11476] = 'b110000010;assign rom[11477] = 'b111000000;assign rom[11478] = 'b101001100;assign rom[11479] = 'b001001010;assign rom[11480] = 'b111111000;assign rom[11481] = 'b111101000;assign rom[11482] = 'b101001111;assign rom[11483] = 'b000111010;assign rom[11484] = 'b101110110;assign rom[11485] = 'b101100010;assign rom[11486] = 'b101001100;assign rom[11487] = 'b001001010;assign rom[11488] = 'b111011010;assign rom[11489] = 'b111011010;assign rom[11490] = 'b111011010;assign rom[11491] = 'b111011010;assign rom[11492] = 'b111011000;assign rom[11493] = 'b111011000;assign rom[11494] = 'b111011000;assign rom[11495] = 'b111011000;assign rom[11496] = 'b101111000;assign rom[11497] = 'b000110011;assign rom[11498] = 'b110000010;assign rom[11499] = 'b001101010;assign rom[11500] = 'b001011000;assign rom[11501] = 'b101001000;assign rom[11502] = 'b000101011;assign rom[11503] = 'b110000010;assign rom[11504] = 'b111000000;assign rom[11505] = 'b101001100;assign rom[11506] = 'b001001010;assign rom[11507] = 'b111111000;assign rom[11508] = 'b111101000;assign rom[11509] = 'b101001111;assign rom[11510] = 'b000111010;assign rom[11511] = 'b101110110;assign rom[11512] = 'b101100010;assign rom[11513] = 'b101001100;assign rom[11514] = 'b001001010;assign rom[11515] = 'b111011010;assign rom[11516] = 'b111011010;assign rom[11517] = 'b111011010;assign rom[11518] = 'b111011010;assign rom[11519] = 'b111011000;assign rom[11520] = 'b111011000;assign rom[11521] = 'b111011000;assign rom[11522] = 'b111011000;assign rom[11523] = 'b101111000;assign rom[11524] = 'b000110011;assign rom[11525] = 'b110000010;assign rom[11526] = 'b001101010;assign rom[11527] = 'b001011000;assign rom[11528] = 'b101001000;assign rom[11529] = 'b000101011;assign rom[11530] = 'b110000010;assign rom[11531] = 'b111000000;assign rom[11532] = 'b101001100;assign rom[11533] = 'b001001010;assign rom[11534] = 'b111111000;assign rom[11535] = 'b111101000;assign rom[11536] = 'b101001111;assign rom[11537] = 'b000111010;assign rom[11538] = 'b101110110;assign rom[11539] = 'b101100010;assign rom[11540] = 'b101001100;assign rom[11541] = 'b001001010;assign rom[11542] = 'b111011010;assign rom[11543] = 'b111011010;assign rom[11544] = 'b111011010;assign rom[11545] = 'b111011010;assign rom[11546] = 'b111011000;assign rom[11547] = 'b111011000;assign rom[11548] = 'b111011000;assign rom[11549] = 'b111011000;assign rom[11550] = 'b101111000;assign rom[11551] = 'b000110011;assign rom[11552] = 'b110000010;assign rom[11553] = 'b001101010;assign rom[11554] = 'b001011000;assign rom[11555] = 'b101001000;assign rom[11556] = 'b000101011;assign rom[11557] = 'b110000010;assign rom[11558] = 'b111000000;assign rom[11559] = 'b101001100;assign rom[11560] = 'b001001010;assign rom[11561] = 'b001000110;assign rom[11562] = 'b001100100;assign rom[11563] = 'b101100010;assign rom[11564] = 'b101001100;assign rom[11565] = 'b001001010;assign rom[11566] = 'b111011010;assign rom[11567] = 'b111011010;assign rom[11568] = 'b111011010;assign rom[11569] = 'b111011010;assign rom[11570] = 'b111011000;assign rom[11571] = 'b111011000;assign rom[11572] = 'b111011000;assign rom[11573] = 'b111011000;assign rom[11574] = 'b101111000;assign rom[11575] = 'b000110011;assign rom[11576] = 'b110000010;assign rom[11577] = 'b001101010;assign rom[11578] = 'b001011000;assign rom[11579] = 'b101001000;assign rom[11580] = 'b000101011;assign rom[11581] = 'b110000010;assign rom[11582] = 'b111000000;assign rom[11583] = 'b101001100;assign rom[11584] = 'b001001010;assign rom[11585] = 'b111111000;assign rom[11586] = 'b111101000;assign rom[11587] = 'b101001111;assign rom[11588] = 'b000111010;assign rom[11589] = 'b101110110;assign rom[11590] = 'b101100010;assign rom[11591] = 'b101001100;assign rom[11592] = 'b001001010;assign rom[11593] = 'b111011010;assign rom[11594] = 'b111011010;assign rom[11595] = 'b111011010;assign rom[11596] = 'b111011010;assign rom[11597] = 'b111011000;assign rom[11598] = 'b111011000;assign rom[11599] = 'b111011000;assign rom[11600] = 'b111011000;assign rom[11601] = 'b101111000;assign rom[11602] = 'b000110011;assign rom[11603] = 'b110000010;assign rom[11604] = 'b001101010;assign rom[11605] = 'b001011000;assign rom[11606] = 'b101001000;assign rom[11607] = 'b000101011;assign rom[11608] = 'b110000010;assign rom[11609] = 'b111000000;assign rom[11610] = 'b101001100;assign rom[11611] = 'b001001010;assign rom[11612] = 'b111111000;assign rom[11613] = 'b111101000;assign rom[11614] = 'b101001111;assign rom[11615] = 'b000111010;assign rom[11616] = 'b101110110;assign rom[11617] = 'b101100010;assign rom[11618] = 'b101001100;assign rom[11619] = 'b001001010;assign rom[11620] = 'b111011010;assign rom[11621] = 'b111011010;assign rom[11622] = 'b111011010;assign rom[11623] = 'b111011010;assign rom[11624] = 'b111011000;assign rom[11625] = 'b111011000;assign rom[11626] = 'b111011000;assign rom[11627] = 'b111011000;assign rom[11628] = 'b101111000;assign rom[11629] = 'b000110011;assign rom[11630] = 'b110000010;assign rom[11631] = 'b001101010;assign rom[11632] = 'b001011000;assign rom[11633] = 'b101001000;assign rom[11634] = 'b000101011;assign rom[11635] = 'b110000010;assign rom[11636] = 'b111000000;assign rom[11637] = 'b101001100;assign rom[11638] = 'b001001010;assign rom[11639] = 'b111111000;assign rom[11640] = 'b111101000;assign rom[11641] = 'b101001111;assign rom[11642] = 'b000111010;assign rom[11643] = 'b101110110;assign rom[11644] = 'b101100010;assign rom[11645] = 'b101001100;assign rom[11646] = 'b001001010;assign rom[11647] = 'b111011010;assign rom[11648] = 'b111011010;assign rom[11649] = 'b111011010;assign rom[11650] = 'b111011010;assign rom[11651] = 'b111011000;assign rom[11652] = 'b111011000;assign rom[11653] = 'b111011000;assign rom[11654] = 'b111011000;assign rom[11655] = 'b101111000;assign rom[11656] = 'b000110011;assign rom[11657] = 'b110000010;assign rom[11658] = 'b001101010;assign rom[11659] = 'b001011000;assign rom[11660] = 'b101001000;assign rom[11661] = 'b000101011;assign rom[11662] = 'b110000010;assign rom[11663] = 'b111000000;assign rom[11664] = 'b101001100;assign rom[11665] = 'b001001010;assign rom[11666] = 'b111111000;assign rom[11667] = 'b111101000;assign rom[11668] = 'b101001111;assign rom[11669] = 'b000111010;assign rom[11670] = 'b101110110;assign rom[11671] = 'b101100010;assign rom[11672] = 'b101001100;assign rom[11673] = 'b001001010;assign rom[11674] = 'b111011010;assign rom[11675] = 'b111011010;assign rom[11676] = 'b111011010;assign rom[11677] = 'b111011010;assign rom[11678] = 'b111011000;assign rom[11679] = 'b111011000;assign rom[11680] = 'b111011000;assign rom[11681] = 'b111011000;assign rom[11682] = 'b101111000;assign rom[11683] = 'b000110011;assign rom[11684] = 'b110000010;assign rom[11685] = 'b001101010;assign rom[11686] = 'b001011000;assign rom[11687] = 'b101001000;assign rom[11688] = 'b000101011;assign rom[11689] = 'b110000010;assign rom[11690] = 'b111000000;assign rom[11691] = 'b101001100;assign rom[11692] = 'b001001010;assign rom[11693] = 'b111111000;assign rom[11694] = 'b111101000;assign rom[11695] = 'b101001111;assign rom[11696] = 'b000111010;assign rom[11697] = 'b101110110;assign rom[11698] = 'b101100010;assign rom[11699] = 'b101001100;assign rom[11700] = 'b001001010;assign rom[11701] = 'b111011010;assign rom[11702] = 'b111011010;assign rom[11703] = 'b111011010;assign rom[11704] = 'b111011010;assign rom[11705] = 'b111011000;assign rom[11706] = 'b111011000;assign rom[11707] = 'b111011000;assign rom[11708] = 'b111011000;assign rom[11709] = 'b101111000;assign rom[11710] = 'b000110011;assign rom[11711] = 'b110000010;assign rom[11712] = 'b001101010;assign rom[11713] = 'b001011000;assign rom[11714] = 'b101001000;assign rom[11715] = 'b000101011;assign rom[11716] = 'b110000010;assign rom[11717] = 'b111000000;assign rom[11718] = 'b101001100;assign rom[11719] = 'b001001010;assign rom[11720] = 'b111111000;assign rom[11721] = 'b111101000;assign rom[11722] = 'b101001111;assign rom[11723] = 'b000111010;assign rom[11724] = 'b101110110;assign rom[11725] = 'b101100010;assign rom[11726] = 'b101001100;assign rom[11727] = 'b001001010;assign rom[11728] = 'b111011010;assign rom[11729] = 'b111011010;assign rom[11730] = 'b111011010;assign rom[11731] = 'b111011010;assign rom[11732] = 'b111011000;assign rom[11733] = 'b111011000;assign rom[11734] = 'b111011000;assign rom[11735] = 'b111011000;assign rom[11736] = 'b101111000;assign rom[11737] = 'b000110011;assign rom[11738] = 'b110000010;assign rom[11739] = 'b001101010;assign rom[11740] = 'b001011000;assign rom[11741] = 'b101001000;assign rom[11742] = 'b000101011;assign rom[11743] = 'b110000010;assign rom[11744] = 'b111000000;assign rom[11745] = 'b101001100;assign rom[11746] = 'b001001010;assign rom[11747] = 'b111111000;assign rom[11748] = 'b111101000;assign rom[11749] = 'b101001111;assign rom[11750] = 'b000111010;assign rom[11751] = 'b101110110;assign rom[11752] = 'b101100010;assign rom[11753] = 'b101001100;assign rom[11754] = 'b001001010;assign rom[11755] = 'b111011010;assign rom[11756] = 'b111011010;assign rom[11757] = 'b111011010;assign rom[11758] = 'b111011010;assign rom[11759] = 'b111011000;assign rom[11760] = 'b111011000;assign rom[11761] = 'b111011000;assign rom[11762] = 'b111011000;assign rom[11763] = 'b101111000;assign rom[11764] = 'b000110011;assign rom[11765] = 'b110000010;assign rom[11766] = 'b001101010;assign rom[11767] = 'b001011000;assign rom[11768] = 'b101001000;assign rom[11769] = 'b000101011;assign rom[11770] = 'b110000010;assign rom[11771] = 'b111000000;assign rom[11772] = 'b101001100;assign rom[11773] = 'b001001010;assign rom[11774] = 'b111111000;assign rom[11775] = 'b111101000;assign rom[11776] = 'b101001111;assign rom[11777] = 'b000111010;assign rom[11778] = 'b101110110;assign rom[11779] = 'b101100010;assign rom[11780] = 'b101001100;assign rom[11781] = 'b001001010;assign rom[11782] = 'b111011010;assign rom[11783] = 'b111011010;assign rom[11784] = 'b111011010;assign rom[11785] = 'b111011010;assign rom[11786] = 'b111011000;assign rom[11787] = 'b111011000;assign rom[11788] = 'b111011000;assign rom[11789] = 'b111011000;assign rom[11790] = 'b101111000;assign rom[11791] = 'b000110011;assign rom[11792] = 'b110000010;assign rom[11793] = 'b001101010;assign rom[11794] = 'b001011000;assign rom[11795] = 'b101001000;assign rom[11796] = 'b000101011;assign rom[11797] = 'b110000010;assign rom[11798] = 'b111000000;assign rom[11799] = 'b101001100;assign rom[11800] = 'b001001010;assign rom[11801] = 'b001000110;assign rom[11802] = 'b001100100;assign rom[11803] = 'b101100010;assign rom[11804] = 'b101001100;assign rom[11805] = 'b001001010;assign rom[11806] = 'b111011010;assign rom[11807] = 'b111011010;assign rom[11808] = 'b111011010;assign rom[11809] = 'b111011010;assign rom[11810] = 'b111011000;assign rom[11811] = 'b111011000;assign rom[11812] = 'b111011000;assign rom[11813] = 'b111011000;assign rom[11814] = 'b101111000;assign rom[11815] = 'b000110011;assign rom[11816] = 'b110000010;assign rom[11817] = 'b001101010;assign rom[11818] = 'b001011000;assign rom[11819] = 'b101001000;assign rom[11820] = 'b000101011;assign rom[11821] = 'b110000010;assign rom[11822] = 'b111000000;assign rom[11823] = 'b101001100;assign rom[11824] = 'b001001010;assign rom[11825] = 'b111111000;assign rom[11826] = 'b111101000;assign rom[11827] = 'b101001111;assign rom[11828] = 'b000111010;assign rom[11829] = 'b101110110;assign rom[11830] = 'b101100010;assign rom[11831] = 'b101001100;assign rom[11832] = 'b001001010;assign rom[11833] = 'b111011010;assign rom[11834] = 'b111011010;assign rom[11835] = 'b111011010;assign rom[11836] = 'b111011010;assign rom[11837] = 'b111011000;assign rom[11838] = 'b111011000;assign rom[11839] = 'b111011000;assign rom[11840] = 'b111011000;assign rom[11841] = 'b101111000;assign rom[11842] = 'b000110011;assign rom[11843] = 'b110000010;assign rom[11844] = 'b001101010;assign rom[11845] = 'b001011000;assign rom[11846] = 'b101001000;assign rom[11847] = 'b000101011;assign rom[11848] = 'b110000010;assign rom[11849] = 'b111000000;assign rom[11850] = 'b101001100;assign rom[11851] = 'b001001010;assign rom[11852] = 'b111111000;assign rom[11853] = 'b111101000;assign rom[11854] = 'b101001111;assign rom[11855] = 'b000111010;assign rom[11856] = 'b101110110;assign rom[11857] = 'b101100010;assign rom[11858] = 'b101001100;assign rom[11859] = 'b001001010;assign rom[11860] = 'b111011010;assign rom[11861] = 'b111011010;assign rom[11862] = 'b111011010;assign rom[11863] = 'b111011010;assign rom[11864] = 'b111011000;assign rom[11865] = 'b111011000;assign rom[11866] = 'b111011000;assign rom[11867] = 'b111011000;assign rom[11868] = 'b101111000;assign rom[11869] = 'b000110011;assign rom[11870] = 'b110000010;assign rom[11871] = 'b001101010;assign rom[11872] = 'b001011000;assign rom[11873] = 'b101001000;assign rom[11874] = 'b000101011;assign rom[11875] = 'b110000010;assign rom[11876] = 'b111000000;assign rom[11877] = 'b101001100;assign rom[11878] = 'b001001010;assign rom[11879] = 'b111111000;assign rom[11880] = 'b111101000;assign rom[11881] = 'b101001111;assign rom[11882] = 'b000111010;assign rom[11883] = 'b101110110;assign rom[11884] = 'b101100010;assign rom[11885] = 'b101001100;assign rom[11886] = 'b001001010;assign rom[11887] = 'b111011010;assign rom[11888] = 'b111011010;assign rom[11889] = 'b111011010;assign rom[11890] = 'b111011010;assign rom[11891] = 'b111011000;assign rom[11892] = 'b111011000;assign rom[11893] = 'b111011000;assign rom[11894] = 'b111011000;assign rom[11895] = 'b101111000;assign rom[11896] = 'b000110011;assign rom[11897] = 'b110000010;assign rom[11898] = 'b001101010;assign rom[11899] = 'b001011000;assign rom[11900] = 'b101001000;assign rom[11901] = 'b000101011;assign rom[11902] = 'b110000010;assign rom[11903] = 'b111000000;assign rom[11904] = 'b101001100;assign rom[11905] = 'b001001010;assign rom[11906] = 'b111111000;assign rom[11907] = 'b111101000;assign rom[11908] = 'b101001111;assign rom[11909] = 'b000111010;assign rom[11910] = 'b101110110;assign rom[11911] = 'b101100010;assign rom[11912] = 'b101001100;assign rom[11913] = 'b001001010;assign rom[11914] = 'b111011010;assign rom[11915] = 'b111011010;assign rom[11916] = 'b111011010;assign rom[11917] = 'b111011010;assign rom[11918] = 'b111011000;assign rom[11919] = 'b111011000;assign rom[11920] = 'b111011000;assign rom[11921] = 'b111011000;assign rom[11922] = 'b101111000;assign rom[11923] = 'b000110011;assign rom[11924] = 'b110000010;assign rom[11925] = 'b001101010;assign rom[11926] = 'b001011000;assign rom[11927] = 'b101001000;assign rom[11928] = 'b000101011;assign rom[11929] = 'b110000010;assign rom[11930] = 'b111000000;assign rom[11931] = 'b101001100;assign rom[11932] = 'b001001010;assign rom[11933] = 'b111111000;assign rom[11934] = 'b111101000;assign rom[11935] = 'b101001111;assign rom[11936] = 'b000111010;assign rom[11937] = 'b101110110;assign rom[11938] = 'b101100010;assign rom[11939] = 'b101001100;assign rom[11940] = 'b001001010;assign rom[11941] = 'b111011010;assign rom[11942] = 'b111011010;assign rom[11943] = 'b111011010;assign rom[11944] = 'b111011010;assign rom[11945] = 'b111011000;assign rom[11946] = 'b111011000;assign rom[11947] = 'b111011000;assign rom[11948] = 'b111011000;assign rom[11949] = 'b101111000;assign rom[11950] = 'b000110011;assign rom[11951] = 'b110000010;assign rom[11952] = 'b001101010;assign rom[11953] = 'b001011000;assign rom[11954] = 'b101001000;assign rom[11955] = 'b000101011;assign rom[11956] = 'b110000010;assign rom[11957] = 'b111000000;assign rom[11958] = 'b101001100;assign rom[11959] = 'b001001010;assign rom[11960] = 'b111111000;assign rom[11961] = 'b111101000;assign rom[11962] = 'b101001111;assign rom[11963] = 'b000111010;assign rom[11964] = 'b101110110;assign rom[11965] = 'b101100010;assign rom[11966] = 'b101001100;assign rom[11967] = 'b001001010;assign rom[11968] = 'b111011010;assign rom[11969] = 'b111011010;assign rom[11970] = 'b111011010;assign rom[11971] = 'b111011010;assign rom[11972] = 'b111011000;assign rom[11973] = 'b111011000;assign rom[11974] = 'b111011000;assign rom[11975] = 'b111011000;assign rom[11976] = 'b101111000;assign rom[11977] = 'b000110011;assign rom[11978] = 'b110000010;assign rom[11979] = 'b001101010;assign rom[11980] = 'b001011000;assign rom[11981] = 'b101001000;assign rom[11982] = 'b000101011;assign rom[11983] = 'b110000010;assign rom[11984] = 'b111000000;assign rom[11985] = 'b101001100;assign rom[11986] = 'b001001010;assign rom[11987] = 'b111111000;assign rom[11988] = 'b111101000;assign rom[11989] = 'b101001111;assign rom[11990] = 'b000111010;assign rom[11991] = 'b101110110;assign rom[11992] = 'b101100010;assign rom[11993] = 'b101001100;assign rom[11994] = 'b001001010;assign rom[11995] = 'b111011010;assign rom[11996] = 'b111011010;assign rom[11997] = 'b111011010;assign rom[11998] = 'b111011010;assign rom[11999] = 'b111011000;assign rom[12000] = 'b111011000;assign rom[12001] = 'b111011000;assign rom[12002] = 'b111011000;assign rom[12003] = 'b101111000;assign rom[12004] = 'b000110011;assign rom[12005] = 'b110000010;assign rom[12006] = 'b001101010;assign rom[12007] = 'b001011000;assign rom[12008] = 'b101001000;assign rom[12009] = 'b000101011;assign rom[12010] = 'b110000010;assign rom[12011] = 'b111000000;assign rom[12012] = 'b101001100;assign rom[12013] = 'b001001010;assign rom[12014] = 'b111111000;assign rom[12015] = 'b111101000;assign rom[12016] = 'b101001111;assign rom[12017] = 'b000111010;assign rom[12018] = 'b101110110;assign rom[12019] = 'b101100010;assign rom[12020] = 'b101001100;assign rom[12021] = 'b001001010;assign rom[12022] = 'b111011010;assign rom[12023] = 'b111011010;assign rom[12024] = 'b111011010;assign rom[12025] = 'b111011010;assign rom[12026] = 'b111011000;assign rom[12027] = 'b111011000;assign rom[12028] = 'b111011000;assign rom[12029] = 'b111011000;assign rom[12030] = 'b101111000;assign rom[12031] = 'b000110011;assign rom[12032] = 'b110000010;assign rom[12033] = 'b001101010;assign rom[12034] = 'b001011000;assign rom[12035] = 'b101001000;assign rom[12036] = 'b000101011;assign rom[12037] = 'b110000010;assign rom[12038] = 'b111000000;assign rom[12039] = 'b101001100;assign rom[12040] = 'b001001010;assign rom[12041] = 'b001000110;assign rom[12042] = 'b001100100;assign rom[12043] = 'b101100010;assign rom[12044] = 'b101001100;assign rom[12045] = 'b001001010;assign rom[12046] = 'b111011010;assign rom[12047] = 'b111011010;assign rom[12048] = 'b111011010;assign rom[12049] = 'b111011010;assign rom[12050] = 'b111011000;assign rom[12051] = 'b111011000;assign rom[12052] = 'b111011000;assign rom[12053] = 'b111011000;assign rom[12054] = 'b101111000;assign rom[12055] = 'b000110011;assign rom[12056] = 'b110000010;assign rom[12057] = 'b001101010;assign rom[12058] = 'b001011000;assign rom[12059] = 'b101001000;assign rom[12060] = 'b000101011;assign rom[12061] = 'b110000010;assign rom[12062] = 'b111000000;assign rom[12063] = 'b101001100;assign rom[12064] = 'b001001010;assign rom[12065] = 'b111111000;assign rom[12066] = 'b111101000;assign rom[12067] = 'b101001111;assign rom[12068] = 'b000111010;assign rom[12069] = 'b101110110;assign rom[12070] = 'b101100010;assign rom[12071] = 'b101001100;assign rom[12072] = 'b001001010;assign rom[12073] = 'b111011010;assign rom[12074] = 'b111011010;assign rom[12075] = 'b111011010;assign rom[12076] = 'b111011010;assign rom[12077] = 'b111011000;assign rom[12078] = 'b111011000;assign rom[12079] = 'b111011000;assign rom[12080] = 'b111011000;assign rom[12081] = 'b101111000;assign rom[12082] = 'b000110011;assign rom[12083] = 'b110000010;assign rom[12084] = 'b001101010;assign rom[12085] = 'b001011000;assign rom[12086] = 'b101001000;assign rom[12087] = 'b000101011;assign rom[12088] = 'b110000010;assign rom[12089] = 'b111000000;assign rom[12090] = 'b101001100;assign rom[12091] = 'b001001010;assign rom[12092] = 'b111111000;assign rom[12093] = 'b111101000;assign rom[12094] = 'b101001111;assign rom[12095] = 'b000111010;assign rom[12096] = 'b101110110;assign rom[12097] = 'b101100010;assign rom[12098] = 'b101001100;assign rom[12099] = 'b001001010;assign rom[12100] = 'b111011010;assign rom[12101] = 'b111011010;assign rom[12102] = 'b111011010;assign rom[12103] = 'b111011010;assign rom[12104] = 'b111011000;assign rom[12105] = 'b111011000;assign rom[12106] = 'b111011000;assign rom[12107] = 'b111011000;assign rom[12108] = 'b101111000;assign rom[12109] = 'b000110011;assign rom[12110] = 'b110000010;assign rom[12111] = 'b001101010;assign rom[12112] = 'b001011000;assign rom[12113] = 'b101001000;assign rom[12114] = 'b000101011;assign rom[12115] = 'b110000010;assign rom[12116] = 'b111000000;assign rom[12117] = 'b101001100;assign rom[12118] = 'b001001010;assign rom[12119] = 'b111111000;assign rom[12120] = 'b111101000;assign rom[12121] = 'b101001111;assign rom[12122] = 'b000111010;assign rom[12123] = 'b101110110;assign rom[12124] = 'b101100010;assign rom[12125] = 'b101001100;assign rom[12126] = 'b001001010;assign rom[12127] = 'b111011010;assign rom[12128] = 'b111011010;assign rom[12129] = 'b111011010;assign rom[12130] = 'b111011010;assign rom[12131] = 'b111011000;assign rom[12132] = 'b111011000;assign rom[12133] = 'b111011000;assign rom[12134] = 'b111011000;assign rom[12135] = 'b101111000;assign rom[12136] = 'b000110011;assign rom[12137] = 'b110000010;assign rom[12138] = 'b001101010;assign rom[12139] = 'b001011000;assign rom[12140] = 'b101001000;assign rom[12141] = 'b000101011;assign rom[12142] = 'b110000010;assign rom[12143] = 'b111000000;assign rom[12144] = 'b101001100;assign rom[12145] = 'b001001010;assign rom[12146] = 'b111111000;assign rom[12147] = 'b111101000;assign rom[12148] = 'b101001111;assign rom[12149] = 'b000111010;assign rom[12150] = 'b101110110;assign rom[12151] = 'b101100010;assign rom[12152] = 'b101001100;assign rom[12153] = 'b001001010;assign rom[12154] = 'b111011010;assign rom[12155] = 'b111011010;assign rom[12156] = 'b111011010;assign rom[12157] = 'b111011010;assign rom[12158] = 'b111011000;assign rom[12159] = 'b111011000;assign rom[12160] = 'b111011000;assign rom[12161] = 'b111011000;assign rom[12162] = 'b101111000;assign rom[12163] = 'b000110011;assign rom[12164] = 'b110000010;assign rom[12165] = 'b001101010;assign rom[12166] = 'b001011000;assign rom[12167] = 'b101001000;assign rom[12168] = 'b000101011;assign rom[12169] = 'b110000010;assign rom[12170] = 'b111000000;assign rom[12171] = 'b101001100;assign rom[12172] = 'b001001010;assign rom[12173] = 'b111111000;assign rom[12174] = 'b111101000;assign rom[12175] = 'b101001111;assign rom[12176] = 'b000111010;assign rom[12177] = 'b101110110;assign rom[12178] = 'b101100010;assign rom[12179] = 'b101001100;assign rom[12180] = 'b001001010;assign rom[12181] = 'b111011010;assign rom[12182] = 'b111011010;assign rom[12183] = 'b111011010;assign rom[12184] = 'b111011010;assign rom[12185] = 'b111011000;assign rom[12186] = 'b111011000;assign rom[12187] = 'b111011000;assign rom[12188] = 'b111011000;assign rom[12189] = 'b101111000;assign rom[12190] = 'b000110011;assign rom[12191] = 'b110000010;assign rom[12192] = 'b001101010;assign rom[12193] = 'b001011000;assign rom[12194] = 'b101001000;assign rom[12195] = 'b000101011;assign rom[12196] = 'b110000010;assign rom[12197] = 'b111000000;assign rom[12198] = 'b101001100;assign rom[12199] = 'b001001010;assign rom[12200] = 'b111111000;assign rom[12201] = 'b111101000;assign rom[12202] = 'b101001111;assign rom[12203] = 'b000111010;assign rom[12204] = 'b101110110;assign rom[12205] = 'b101100010;assign rom[12206] = 'b101001100;assign rom[12207] = 'b001001010;assign rom[12208] = 'b111011010;assign rom[12209] = 'b111011010;assign rom[12210] = 'b111011010;assign rom[12211] = 'b111011010;assign rom[12212] = 'b111011000;assign rom[12213] = 'b111011000;assign rom[12214] = 'b111011000;assign rom[12215] = 'b111011000;assign rom[12216] = 'b101111000;assign rom[12217] = 'b000110011;assign rom[12218] = 'b110000010;assign rom[12219] = 'b001101010;assign rom[12220] = 'b001011000;assign rom[12221] = 'b101001000;assign rom[12222] = 'b000101011;assign rom[12223] = 'b110000010;assign rom[12224] = 'b111000000;assign rom[12225] = 'b101001100;assign rom[12226] = 'b001001010;assign rom[12227] = 'b111111000;assign rom[12228] = 'b111101000;assign rom[12229] = 'b101001111;assign rom[12230] = 'b000111010;assign rom[12231] = 'b101110110;assign rom[12232] = 'b101100010;assign rom[12233] = 'b101001100;assign rom[12234] = 'b001001010;assign rom[12235] = 'b111011010;assign rom[12236] = 'b111011010;assign rom[12237] = 'b111011010;assign rom[12238] = 'b111011010;assign rom[12239] = 'b111011000;assign rom[12240] = 'b111011000;assign rom[12241] = 'b111011000;assign rom[12242] = 'b111011000;assign rom[12243] = 'b101111000;assign rom[12244] = 'b000110011;assign rom[12245] = 'b110000010;assign rom[12246] = 'b001101010;assign rom[12247] = 'b001011000;assign rom[12248] = 'b101001000;assign rom[12249] = 'b000101011;assign rom[12250] = 'b110000010;assign rom[12251] = 'b111000000;assign rom[12252] = 'b101001100;assign rom[12253] = 'b001001010;assign rom[12254] = 'b111111000;assign rom[12255] = 'b111101000;assign rom[12256] = 'b101001111;assign rom[12257] = 'b000111010;assign rom[12258] = 'b101110110;assign rom[12259] = 'b101100010;assign rom[12260] = 'b101001100;assign rom[12261] = 'b001001010;assign rom[12262] = 'b111011010;assign rom[12263] = 'b111011010;assign rom[12264] = 'b111011010;assign rom[12265] = 'b111011010;assign rom[12266] = 'b111011000;assign rom[12267] = 'b111011000;assign rom[12268] = 'b111011000;assign rom[12269] = 'b111011000;assign rom[12270] = 'b101111000;assign rom[12271] = 'b000110011;assign rom[12272] = 'b110000010;assign rom[12273] = 'b001101010;assign rom[12274] = 'b001011000;assign rom[12275] = 'b101001000;assign rom[12276] = 'b000101011;assign rom[12277] = 'b110000010;assign rom[12278] = 'b111000000;assign rom[12279] = 'b101001100;assign rom[12280] = 'b001001010;assign rom[12281] = 'b001000110;assign rom[12282] = 'b001100100;assign rom[12283] = 'b101100010;assign rom[12284] = 'b101001100;assign rom[12285] = 'b001001010;assign rom[12286] = 'b111011010;assign rom[12287] = 'b111011010;assign rom[12288] = 'b111011010;assign rom[12289] = 'b111011010;assign rom[12290] = 'b111011000;assign rom[12291] = 'b111011000;assign rom[12292] = 'b111011000;assign rom[12293] = 'b111011000;assign rom[12294] = 'b101111000;assign rom[12295] = 'b000110011;assign rom[12296] = 'b110000010;assign rom[12297] = 'b001101010;assign rom[12298] = 'b001011000;assign rom[12299] = 'b101001000;assign rom[12300] = 'b000101011;assign rom[12301] = 'b110000010;assign rom[12302] = 'b111000000;assign rom[12303] = 'b101001100;assign rom[12304] = 'b001001010;assign rom[12305] = 'b111111000;assign rom[12306] = 'b111101000;assign rom[12307] = 'b101001111;assign rom[12308] = 'b000111010;assign rom[12309] = 'b101110110;assign rom[12310] = 'b101100010;assign rom[12311] = 'b101001100;assign rom[12312] = 'b001001010;assign rom[12313] = 'b111011010;assign rom[12314] = 'b111011010;assign rom[12315] = 'b111011010;assign rom[12316] = 'b111011010;assign rom[12317] = 'b111011000;assign rom[12318] = 'b111011000;assign rom[12319] = 'b111011000;assign rom[12320] = 'b111011000;assign rom[12321] = 'b101111000;assign rom[12322] = 'b000110011;assign rom[12323] = 'b110000010;assign rom[12324] = 'b001101010;assign rom[12325] = 'b001011000;assign rom[12326] = 'b101001000;assign rom[12327] = 'b000101011;assign rom[12328] = 'b110000010;assign rom[12329] = 'b111000000;assign rom[12330] = 'b101001100;assign rom[12331] = 'b001001010;assign rom[12332] = 'b111111000;assign rom[12333] = 'b111101000;assign rom[12334] = 'b101001111;assign rom[12335] = 'b000111010;assign rom[12336] = 'b101110110;assign rom[12337] = 'b101100010;assign rom[12338] = 'b101001100;assign rom[12339] = 'b001001010;assign rom[12340] = 'b111011010;assign rom[12341] = 'b111011010;assign rom[12342] = 'b111011010;assign rom[12343] = 'b111011010;assign rom[12344] = 'b111011000;assign rom[12345] = 'b111011000;assign rom[12346] = 'b111011000;assign rom[12347] = 'b111011000;assign rom[12348] = 'b101111000;assign rom[12349] = 'b000110011;assign rom[12350] = 'b110000010;assign rom[12351] = 'b001101010;assign rom[12352] = 'b001011000;assign rom[12353] = 'b101001000;assign rom[12354] = 'b000101011;assign rom[12355] = 'b110000010;assign rom[12356] = 'b111000000;assign rom[12357] = 'b101001100;assign rom[12358] = 'b001001010;assign rom[12359] = 'b111111000;assign rom[12360] = 'b111101000;assign rom[12361] = 'b101001111;assign rom[12362] = 'b000111010;assign rom[12363] = 'b101110110;assign rom[12364] = 'b101100010;assign rom[12365] = 'b101001100;assign rom[12366] = 'b001001010;assign rom[12367] = 'b111011010;assign rom[12368] = 'b111011010;assign rom[12369] = 'b111011010;assign rom[12370] = 'b111011010;assign rom[12371] = 'b111011000;assign rom[12372] = 'b111011000;assign rom[12373] = 'b111011000;assign rom[12374] = 'b111011000;assign rom[12375] = 'b101111000;assign rom[12376] = 'b000110011;assign rom[12377] = 'b110000010;assign rom[12378] = 'b001101010;assign rom[12379] = 'b001011000;assign rom[12380] = 'b101001000;assign rom[12381] = 'b000101011;assign rom[12382] = 'b110000010;assign rom[12383] = 'b111000000;assign rom[12384] = 'b101001100;assign rom[12385] = 'b001001010;assign rom[12386] = 'b111111000;assign rom[12387] = 'b111101000;assign rom[12388] = 'b101001111;assign rom[12389] = 'b000111010;assign rom[12390] = 'b101110110;assign rom[12391] = 'b101100010;assign rom[12392] = 'b101001100;assign rom[12393] = 'b001001010;assign rom[12394] = 'b111011010;assign rom[12395] = 'b111011010;assign rom[12396] = 'b111011010;assign rom[12397] = 'b111011010;assign rom[12398] = 'b111011000;assign rom[12399] = 'b111011000;assign rom[12400] = 'b111011000;assign rom[12401] = 'b111011000;assign rom[12402] = 'b101111000;assign rom[12403] = 'b000110011;assign rom[12404] = 'b110000010;assign rom[12405] = 'b001101010;assign rom[12406] = 'b001011000;assign rom[12407] = 'b101001000;assign rom[12408] = 'b000101011;assign rom[12409] = 'b110000010;assign rom[12410] = 'b111000000;assign rom[12411] = 'b101001100;assign rom[12412] = 'b001001010;assign rom[12413] = 'b111111000;assign rom[12414] = 'b111101000;assign rom[12415] = 'b101001111;assign rom[12416] = 'b000111010;assign rom[12417] = 'b101110110;assign rom[12418] = 'b101100010;assign rom[12419] = 'b101001100;assign rom[12420] = 'b001001010;assign rom[12421] = 'b111011010;assign rom[12422] = 'b111011010;assign rom[12423] = 'b111011010;assign rom[12424] = 'b111011010;assign rom[12425] = 'b111011000;assign rom[12426] = 'b111011000;assign rom[12427] = 'b111011000;assign rom[12428] = 'b111011000;assign rom[12429] = 'b101111000;assign rom[12430] = 'b000110011;assign rom[12431] = 'b110000010;assign rom[12432] = 'b001101010;assign rom[12433] = 'b001011000;assign rom[12434] = 'b101001000;assign rom[12435] = 'b000101011;assign rom[12436] = 'b110000010;assign rom[12437] = 'b111000000;assign rom[12438] = 'b101001100;assign rom[12439] = 'b001001010;assign rom[12440] = 'b111111000;assign rom[12441] = 'b111101000;assign rom[12442] = 'b101001111;assign rom[12443] = 'b000111010;assign rom[12444] = 'b101110110;assign rom[12445] = 'b101100010;assign rom[12446] = 'b101001100;assign rom[12447] = 'b001001010;assign rom[12448] = 'b111011010;assign rom[12449] = 'b111011010;assign rom[12450] = 'b111011010;assign rom[12451] = 'b111011010;assign rom[12452] = 'b111011000;assign rom[12453] = 'b111011000;assign rom[12454] = 'b111011000;assign rom[12455] = 'b111011000;assign rom[12456] = 'b101111000;assign rom[12457] = 'b000110011;assign rom[12458] = 'b110000010;assign rom[12459] = 'b001101010;assign rom[12460] = 'b001011000;assign rom[12461] = 'b101001000;assign rom[12462] = 'b000101011;assign rom[12463] = 'b110000010;assign rom[12464] = 'b111000000;assign rom[12465] = 'b101001100;assign rom[12466] = 'b001001010;assign rom[12467] = 'b111111000;assign rom[12468] = 'b111101000;assign rom[12469] = 'b101001111;assign rom[12470] = 'b000111010;assign rom[12471] = 'b101110110;assign rom[12472] = 'b101100010;assign rom[12473] = 'b101001100;assign rom[12474] = 'b001001010;assign rom[12475] = 'b111011010;assign rom[12476] = 'b111011010;assign rom[12477] = 'b111011010;assign rom[12478] = 'b111011010;assign rom[12479] = 'b111011000;assign rom[12480] = 'b111011000;assign rom[12481] = 'b111011000;assign rom[12482] = 'b111011000;assign rom[12483] = 'b101111000;assign rom[12484] = 'b000110011;assign rom[12485] = 'b110000010;assign rom[12486] = 'b001101010;assign rom[12487] = 'b001011000;assign rom[12488] = 'b101001000;assign rom[12489] = 'b000101011;assign rom[12490] = 'b110000010;assign rom[12491] = 'b111000000;assign rom[12492] = 'b101001100;assign rom[12493] = 'b001001010;assign rom[12494] = 'b111111000;assign rom[12495] = 'b111101000;assign rom[12496] = 'b101001111;assign rom[12497] = 'b000111010;assign rom[12498] = 'b101110110;assign rom[12499] = 'b101100010;assign rom[12500] = 'b101001100;assign rom[12501] = 'b001001010;assign rom[12502] = 'b111011010;assign rom[12503] = 'b111011010;assign rom[12504] = 'b111011010;assign rom[12505] = 'b111011010;assign rom[12506] = 'b111011000;assign rom[12507] = 'b111011000;assign rom[12508] = 'b111011000;assign rom[12509] = 'b111011000;assign rom[12510] = 'b101111000;assign rom[12511] = 'b000110011;assign rom[12512] = 'b110000010;assign rom[12513] = 'b001101010;assign rom[12514] = 'b001011000;assign rom[12515] = 'b101001000;assign rom[12516] = 'b000101011;assign rom[12517] = 'b110000010;assign rom[12518] = 'b111000000;assign rom[12519] = 'b101001100;assign rom[12520] = 'b001001010;assign rom[12521] = 'b001000110;assign rom[12522] = 'b001100100;assign rom[12523] = 'b101100010;assign rom[12524] = 'b101001100;assign rom[12525] = 'b001001010;assign rom[12526] = 'b111011010;assign rom[12527] = 'b111011010;assign rom[12528] = 'b111011010;assign rom[12529] = 'b111011010;assign rom[12530] = 'b111011000;assign rom[12531] = 'b111011000;assign rom[12532] = 'b111011000;assign rom[12533] = 'b111011000;assign rom[12534] = 'b101111000;assign rom[12535] = 'b000110011;assign rom[12536] = 'b110000010;assign rom[12537] = 'b001101010;assign rom[12538] = 'b001011000;assign rom[12539] = 'b101001000;assign rom[12540] = 'b000101011;assign rom[12541] = 'b110000010;assign rom[12542] = 'b111000000;assign rom[12543] = 'b101001100;assign rom[12544] = 'b001001010;assign rom[12545] = 'b111111000;assign rom[12546] = 'b111101000;assign rom[12547] = 'b101001111;assign rom[12548] = 'b000111010;assign rom[12549] = 'b101110110;assign rom[12550] = 'b101100010;assign rom[12551] = 'b101001100;assign rom[12552] = 'b001001010;assign rom[12553] = 'b111011010;assign rom[12554] = 'b111011010;assign rom[12555] = 'b111011010;assign rom[12556] = 'b111011010;assign rom[12557] = 'b111011000;assign rom[12558] = 'b111011000;assign rom[12559] = 'b111011000;assign rom[12560] = 'b111011000;assign rom[12561] = 'b101111000;assign rom[12562] = 'b000110011;assign rom[12563] = 'b110000010;assign rom[12564] = 'b001101010;assign rom[12565] = 'b001011000;assign rom[12566] = 'b101001000;assign rom[12567] = 'b000101011;assign rom[12568] = 'b110000010;assign rom[12569] = 'b111000000;assign rom[12570] = 'b101001100;assign rom[12571] = 'b001001010;assign rom[12572] = 'b111111000;assign rom[12573] = 'b111101000;assign rom[12574] = 'b101001111;assign rom[12575] = 'b000111010;assign rom[12576] = 'b101110110;assign rom[12577] = 'b101100010;assign rom[12578] = 'b101001100;assign rom[12579] = 'b001001010;assign rom[12580] = 'b111011010;assign rom[12581] = 'b111011010;assign rom[12582] = 'b111011010;assign rom[12583] = 'b111011010;assign rom[12584] = 'b111011000;assign rom[12585] = 'b111011000;assign rom[12586] = 'b111011000;assign rom[12587] = 'b111011000;assign rom[12588] = 'b101111000;assign rom[12589] = 'b000110011;assign rom[12590] = 'b110000010;assign rom[12591] = 'b001101010;assign rom[12592] = 'b001011000;assign rom[12593] = 'b101001000;assign rom[12594] = 'b000101011;assign rom[12595] = 'b110000010;assign rom[12596] = 'b111000000;assign rom[12597] = 'b101001100;assign rom[12598] = 'b001001010;assign rom[12599] = 'b111111000;assign rom[12600] = 'b111101000;assign rom[12601] = 'b101001111;assign rom[12602] = 'b000111010;assign rom[12603] = 'b101110110;assign rom[12604] = 'b101100010;assign rom[12605] = 'b101001100;assign rom[12606] = 'b001001010;assign rom[12607] = 'b111011010;assign rom[12608] = 'b111011010;assign rom[12609] = 'b111011010;assign rom[12610] = 'b111011010;assign rom[12611] = 'b111011000;assign rom[12612] = 'b111011000;assign rom[12613] = 'b111011000;assign rom[12614] = 'b111011000;assign rom[12615] = 'b101111000;assign rom[12616] = 'b000110011;assign rom[12617] = 'b110000010;assign rom[12618] = 'b001101010;assign rom[12619] = 'b001011000;assign rom[12620] = 'b101001000;assign rom[12621] = 'b000101011;assign rom[12622] = 'b110000010;assign rom[12623] = 'b111000000;assign rom[12624] = 'b101001100;assign rom[12625] = 'b001001010;assign rom[12626] = 'b111111000;assign rom[12627] = 'b111101000;assign rom[12628] = 'b101001111;assign rom[12629] = 'b000111010;assign rom[12630] = 'b101110110;assign rom[12631] = 'b101100010;assign rom[12632] = 'b101001100;assign rom[12633] = 'b001001010;assign rom[12634] = 'b111011010;assign rom[12635] = 'b111011010;assign rom[12636] = 'b111011010;assign rom[12637] = 'b111011010;assign rom[12638] = 'b111011000;assign rom[12639] = 'b111011000;assign rom[12640] = 'b111011000;assign rom[12641] = 'b111011000;assign rom[12642] = 'b101111000;assign rom[12643] = 'b000110011;assign rom[12644] = 'b110000010;assign rom[12645] = 'b001101010;assign rom[12646] = 'b001011000;assign rom[12647] = 'b101001000;assign rom[12648] = 'b000101011;assign rom[12649] = 'b110000010;assign rom[12650] = 'b111000000;assign rom[12651] = 'b101001100;assign rom[12652] = 'b001001010;assign rom[12653] = 'b111111000;assign rom[12654] = 'b111101000;assign rom[12655] = 'b101001111;assign rom[12656] = 'b000111010;assign rom[12657] = 'b101110110;assign rom[12658] = 'b101100010;assign rom[12659] = 'b101001100;assign rom[12660] = 'b001001010;assign rom[12661] = 'b111011010;assign rom[12662] = 'b111011010;assign rom[12663] = 'b111011010;assign rom[12664] = 'b111011010;assign rom[12665] = 'b111011000;assign rom[12666] = 'b111011000;assign rom[12667] = 'b111011000;assign rom[12668] = 'b111011000;assign rom[12669] = 'b101111000;assign rom[12670] = 'b000110011;assign rom[12671] = 'b110000010;assign rom[12672] = 'b001101010;assign rom[12673] = 'b001011000;assign rom[12674] = 'b101001000;assign rom[12675] = 'b000101011;assign rom[12676] = 'b110000010;assign rom[12677] = 'b111000000;assign rom[12678] = 'b101001100;assign rom[12679] = 'b001001010;assign rom[12680] = 'b111111000;assign rom[12681] = 'b111101000;assign rom[12682] = 'b101001111;assign rom[12683] = 'b000111010;assign rom[12684] = 'b101110110;assign rom[12685] = 'b101100010;assign rom[12686] = 'b101001100;assign rom[12687] = 'b001001010;assign rom[12688] = 'b111011010;assign rom[12689] = 'b111011010;assign rom[12690] = 'b111011010;assign rom[12691] = 'b111011010;assign rom[12692] = 'b111011000;assign rom[12693] = 'b111011000;assign rom[12694] = 'b111011000;assign rom[12695] = 'b111011000;assign rom[12696] = 'b101111000;assign rom[12697] = 'b000110011;assign rom[12698] = 'b110000010;assign rom[12699] = 'b001101010;assign rom[12700] = 'b001011000;assign rom[12701] = 'b101001000;assign rom[12702] = 'b000101011;assign rom[12703] = 'b110000010;assign rom[12704] = 'b111000000;assign rom[12705] = 'b101001100;assign rom[12706] = 'b001001010;assign rom[12707] = 'b111111000;assign rom[12708] = 'b111101000;assign rom[12709] = 'b101001111;assign rom[12710] = 'b000111010;assign rom[12711] = 'b101110110;assign rom[12712] = 'b101100010;assign rom[12713] = 'b101001100;assign rom[12714] = 'b001001010;assign rom[12715] = 'b111011010;assign rom[12716] = 'b111011010;assign rom[12717] = 'b111011010;assign rom[12718] = 'b111011010;assign rom[12719] = 'b111011000;assign rom[12720] = 'b111011000;assign rom[12721] = 'b111011000;assign rom[12722] = 'b111011000;assign rom[12723] = 'b101111000;assign rom[12724] = 'b000110011;assign rom[12725] = 'b110000010;assign rom[12726] = 'b001101010;assign rom[12727] = 'b001011000;assign rom[12728] = 'b101001000;assign rom[12729] = 'b000101011;assign rom[12730] = 'b110000010;assign rom[12731] = 'b111000000;assign rom[12732] = 'b101001100;assign rom[12733] = 'b001001010;assign rom[12734] = 'b111111000;assign rom[12735] = 'b111101000;assign rom[12736] = 'b101001111;assign rom[12737] = 'b000111010;assign rom[12738] = 'b101110110;assign rom[12739] = 'b101100010;assign rom[12740] = 'b101001100;assign rom[12741] = 'b001001010;assign rom[12742] = 'b111011010;assign rom[12743] = 'b111011010;assign rom[12744] = 'b111011010;assign rom[12745] = 'b111011010;assign rom[12746] = 'b111011000;assign rom[12747] = 'b111011000;assign rom[12748] = 'b111011000;assign rom[12749] = 'b111011000;assign rom[12750] = 'b101111000;assign rom[12751] = 'b000110011;assign rom[12752] = 'b110000010;assign rom[12753] = 'b001101010;assign rom[12754] = 'b001011000;assign rom[12755] = 'b101001000;assign rom[12756] = 'b000101011;assign rom[12757] = 'b110000010;assign rom[12758] = 'b111000000;assign rom[12759] = 'b101001100;assign rom[12760] = 'b001001010;assign rom[12761] = 'b001000110;assign rom[12762] = 'b001100100;assign rom[12763] = 'b101100010;assign rom[12764] = 'b101001100;assign rom[12765] = 'b001001010;assign rom[12766] = 'b111011010;assign rom[12767] = 'b111011010;assign rom[12768] = 'b111011010;assign rom[12769] = 'b111011010;assign rom[12770] = 'b111011000;assign rom[12771] = 'b111011000;assign rom[12772] = 'b111011000;assign rom[12773] = 'b111011000;assign rom[12774] = 'b101111000;assign rom[12775] = 'b000110011;assign rom[12776] = 'b110000010;assign rom[12777] = 'b001101010;assign rom[12778] = 'b001011000;assign rom[12779] = 'b101001000;assign rom[12780] = 'b000101011;assign rom[12781] = 'b110000010;assign rom[12782] = 'b111000000;assign rom[12783] = 'b101001100;assign rom[12784] = 'b001001010;assign rom[12785] = 'b111111000;assign rom[12786] = 'b111101000;assign rom[12787] = 'b101001111;assign rom[12788] = 'b000111010;assign rom[12789] = 'b101110110;assign rom[12790] = 'b101100010;assign rom[12791] = 'b101001100;assign rom[12792] = 'b001001010;assign rom[12793] = 'b111011010;assign rom[12794] = 'b111011010;assign rom[12795] = 'b111011010;assign rom[12796] = 'b111011010;assign rom[12797] = 'b111011000;assign rom[12798] = 'b111011000;assign rom[12799] = 'b111011000;assign rom[12800] = 'b111011000;assign rom[12801] = 'b101111000;assign rom[12802] = 'b000110011;assign rom[12803] = 'b110000010;assign rom[12804] = 'b001101010;assign rom[12805] = 'b001011000;assign rom[12806] = 'b101001000;assign rom[12807] = 'b000101011;assign rom[12808] = 'b110000010;assign rom[12809] = 'b111000000;assign rom[12810] = 'b101001100;assign rom[12811] = 'b001001010;assign rom[12812] = 'b111111000;assign rom[12813] = 'b111101000;assign rom[12814] = 'b101001111;assign rom[12815] = 'b000111010;assign rom[12816] = 'b101110110;assign rom[12817] = 'b101100010;assign rom[12818] = 'b101001100;assign rom[12819] = 'b001001010;assign rom[12820] = 'b111011010;assign rom[12821] = 'b111011010;assign rom[12822] = 'b111011010;assign rom[12823] = 'b111011010;assign rom[12824] = 'b111011000;assign rom[12825] = 'b111011000;assign rom[12826] = 'b111011000;assign rom[12827] = 'b111011000;assign rom[12828] = 'b101111000;assign rom[12829] = 'b000110011;assign rom[12830] = 'b110000010;assign rom[12831] = 'b001101010;assign rom[12832] = 'b001011000;assign rom[12833] = 'b101001000;assign rom[12834] = 'b000101011;assign rom[12835] = 'b110000010;assign rom[12836] = 'b111000000;assign rom[12837] = 'b101001100;assign rom[12838] = 'b001001010;assign rom[12839] = 'b111111000;assign rom[12840] = 'b111101000;assign rom[12841] = 'b101001111;assign rom[12842] = 'b000111010;assign rom[12843] = 'b101110110;assign rom[12844] = 'b101100010;assign rom[12845] = 'b101001100;assign rom[12846] = 'b001001010;assign rom[12847] = 'b111011010;assign rom[12848] = 'b111011010;assign rom[12849] = 'b111011010;assign rom[12850] = 'b111011010;assign rom[12851] = 'b111011000;assign rom[12852] = 'b111011000;assign rom[12853] = 'b111011000;assign rom[12854] = 'b111011000;assign rom[12855] = 'b101111000;assign rom[12856] = 'b000110011;assign rom[12857] = 'b110000010;assign rom[12858] = 'b001101010;assign rom[12859] = 'b001011000;assign rom[12860] = 'b101001000;assign rom[12861] = 'b000101011;assign rom[12862] = 'b110000010;assign rom[12863] = 'b111000000;assign rom[12864] = 'b101001100;assign rom[12865] = 'b001001010;assign rom[12866] = 'b111111000;assign rom[12867] = 'b111101000;assign rom[12868] = 'b101001111;assign rom[12869] = 'b000111010;assign rom[12870] = 'b101110110;assign rom[12871] = 'b101100010;assign rom[12872] = 'b101001100;assign rom[12873] = 'b001001010;assign rom[12874] = 'b111011010;assign rom[12875] = 'b111011010;assign rom[12876] = 'b111011010;assign rom[12877] = 'b111011010;assign rom[12878] = 'b111011000;assign rom[12879] = 'b111011000;assign rom[12880] = 'b111011000;assign rom[12881] = 'b111011000;assign rom[12882] = 'b101111000;assign rom[12883] = 'b000110011;assign rom[12884] = 'b110000010;assign rom[12885] = 'b001101010;assign rom[12886] = 'b001011000;assign rom[12887] = 'b101001000;assign rom[12888] = 'b000101011;assign rom[12889] = 'b110000010;assign rom[12890] = 'b111000000;assign rom[12891] = 'b101001100;assign rom[12892] = 'b001001010;assign rom[12893] = 'b111111000;assign rom[12894] = 'b111101000;assign rom[12895] = 'b101001111;assign rom[12896] = 'b000111010;assign rom[12897] = 'b101110110;assign rom[12898] = 'b101100010;assign rom[12899] = 'b101001100;assign rom[12900] = 'b001001010;assign rom[12901] = 'b111011010;assign rom[12902] = 'b111011010;assign rom[12903] = 'b111011010;assign rom[12904] = 'b111011010;assign rom[12905] = 'b111011000;assign rom[12906] = 'b111011000;assign rom[12907] = 'b111011000;assign rom[12908] = 'b111011000;assign rom[12909] = 'b101111000;assign rom[12910] = 'b000110011;assign rom[12911] = 'b110000010;assign rom[12912] = 'b001101010;assign rom[12913] = 'b001011000;assign rom[12914] = 'b101001000;assign rom[12915] = 'b000101011;assign rom[12916] = 'b110000010;assign rom[12917] = 'b111000000;assign rom[12918] = 'b101001100;assign rom[12919] = 'b001001010;assign rom[12920] = 'b111111000;assign rom[12921] = 'b111101000;assign rom[12922] = 'b101001111;assign rom[12923] = 'b000111010;assign rom[12924] = 'b101110110;assign rom[12925] = 'b101100010;assign rom[12926] = 'b101001100;assign rom[12927] = 'b001001010;assign rom[12928] = 'b111011010;assign rom[12929] = 'b111011010;assign rom[12930] = 'b111011010;assign rom[12931] = 'b111011010;assign rom[12932] = 'b111011000;assign rom[12933] = 'b111011000;assign rom[12934] = 'b111011000;assign rom[12935] = 'b111011000;assign rom[12936] = 'b101111000;assign rom[12937] = 'b000110011;assign rom[12938] = 'b110000010;assign rom[12939] = 'b001101010;assign rom[12940] = 'b001011000;assign rom[12941] = 'b101001000;assign rom[12942] = 'b000101011;assign rom[12943] = 'b110000010;assign rom[12944] = 'b111000000;assign rom[12945] = 'b101001100;assign rom[12946] = 'b001001010;assign rom[12947] = 'b111111000;assign rom[12948] = 'b111101000;assign rom[12949] = 'b101001111;assign rom[12950] = 'b000111010;assign rom[12951] = 'b101110110;assign rom[12952] = 'b101100010;assign rom[12953] = 'b101001100;assign rom[12954] = 'b001001010;assign rom[12955] = 'b111011010;assign rom[12956] = 'b111011010;assign rom[12957] = 'b111011010;assign rom[12958] = 'b111011010;assign rom[12959] = 'b111011000;assign rom[12960] = 'b111011000;assign rom[12961] = 'b111011000;assign rom[12962] = 'b111011000;assign rom[12963] = 'b101111000;assign rom[12964] = 'b000110011;assign rom[12965] = 'b110000010;assign rom[12966] = 'b001101010;assign rom[12967] = 'b001011000;assign rom[12968] = 'b101001000;assign rom[12969] = 'b000101011;assign rom[12970] = 'b110000010;assign rom[12971] = 'b111000000;assign rom[12972] = 'b101001100;assign rom[12973] = 'b001001010;assign rom[12974] = 'b111111000;assign rom[12975] = 'b111101000;assign rom[12976] = 'b101001111;assign rom[12977] = 'b000111010;assign rom[12978] = 'b101110110;assign rom[12979] = 'b101100010;assign rom[12980] = 'b101001100;assign rom[12981] = 'b001001010;assign rom[12982] = 'b111011010;assign rom[12983] = 'b111011010;assign rom[12984] = 'b111011010;assign rom[12985] = 'b111011010;assign rom[12986] = 'b111011000;assign rom[12987] = 'b111011000;assign rom[12988] = 'b111011000;assign rom[12989] = 'b111011000;assign rom[12990] = 'b101111000;assign rom[12991] = 'b000110011;assign rom[12992] = 'b110000010;assign rom[12993] = 'b001101010;assign rom[12994] = 'b001011000;assign rom[12995] = 'b101001000;assign rom[12996] = 'b000101011;assign rom[12997] = 'b110000010;assign rom[12998] = 'b111000000;assign rom[12999] = 'b101001100;assign rom[13000] = 'b001001010;assign rom[13001] = 'b001000110;assign rom[13002] = 'b001100100;assign rom[13003] = 'b101100010;assign rom[13004] = 'b101001100;assign rom[13005] = 'b001001010;assign rom[13006] = 'b111011010;assign rom[13007] = 'b111011010;assign rom[13008] = 'b111011010;assign rom[13009] = 'b111011010;assign rom[13010] = 'b111011000;assign rom[13011] = 'b111011000;assign rom[13012] = 'b111011000;assign rom[13013] = 'b111011000;assign rom[13014] = 'b101111000;assign rom[13015] = 'b000110011;assign rom[13016] = 'b110000010;assign rom[13017] = 'b001101010;assign rom[13018] = 'b001011000;assign rom[13019] = 'b101001000;assign rom[13020] = 'b000101011;assign rom[13021] = 'b110000010;assign rom[13022] = 'b111000000;assign rom[13023] = 'b101001100;assign rom[13024] = 'b001001010;assign rom[13025] = 'b111111000;assign rom[13026] = 'b111101000;assign rom[13027] = 'b101001111;assign rom[13028] = 'b000111010;assign rom[13029] = 'b101110110;assign rom[13030] = 'b101100010;assign rom[13031] = 'b101001100;assign rom[13032] = 'b001001010;assign rom[13033] = 'b111011010;assign rom[13034] = 'b111011010;assign rom[13035] = 'b111011010;assign rom[13036] = 'b111011010;assign rom[13037] = 'b111011000;assign rom[13038] = 'b111011000;assign rom[13039] = 'b111011000;assign rom[13040] = 'b111011000;assign rom[13041] = 'b101111000;assign rom[13042] = 'b000110011;assign rom[13043] = 'b110000010;assign rom[13044] = 'b001101010;assign rom[13045] = 'b001011000;assign rom[13046] = 'b101001000;assign rom[13047] = 'b000101011;assign rom[13048] = 'b110000010;assign rom[13049] = 'b111000000;assign rom[13050] = 'b101001100;assign rom[13051] = 'b001001010;assign rom[13052] = 'b111111000;assign rom[13053] = 'b111101000;assign rom[13054] = 'b101001111;assign rom[13055] = 'b000111010;assign rom[13056] = 'b101110110;assign rom[13057] = 'b101100010;assign rom[13058] = 'b101001100;assign rom[13059] = 'b001001010;assign rom[13060] = 'b111011010;assign rom[13061] = 'b111011010;assign rom[13062] = 'b111011010;assign rom[13063] = 'b111011010;assign rom[13064] = 'b111011000;assign rom[13065] = 'b111011000;assign rom[13066] = 'b111011000;assign rom[13067] = 'b111011000;assign rom[13068] = 'b101111000;assign rom[13069] = 'b000110011;assign rom[13070] = 'b110000010;assign rom[13071] = 'b001101010;assign rom[13072] = 'b001011000;assign rom[13073] = 'b101001000;assign rom[13074] = 'b000101011;assign rom[13075] = 'b110000010;assign rom[13076] = 'b111000000;assign rom[13077] = 'b101001100;assign rom[13078] = 'b001001010;assign rom[13079] = 'b111111000;assign rom[13080] = 'b111101000;assign rom[13081] = 'b101001111;assign rom[13082] = 'b000111010;assign rom[13083] = 'b101110110;assign rom[13084] = 'b101100010;assign rom[13085] = 'b101001100;assign rom[13086] = 'b001001010;assign rom[13087] = 'b111011010;assign rom[13088] = 'b111011010;assign rom[13089] = 'b111011010;assign rom[13090] = 'b111011010;assign rom[13091] = 'b111011000;assign rom[13092] = 'b111011000;assign rom[13093] = 'b111011000;assign rom[13094] = 'b111011000;assign rom[13095] = 'b101111000;assign rom[13096] = 'b000110011;assign rom[13097] = 'b110000010;assign rom[13098] = 'b001101010;assign rom[13099] = 'b001011000;assign rom[13100] = 'b101001000;assign rom[13101] = 'b000101011;assign rom[13102] = 'b110000010;assign rom[13103] = 'b111000000;assign rom[13104] = 'b101001100;assign rom[13105] = 'b001001010;assign rom[13106] = 'b111111000;assign rom[13107] = 'b111101000;assign rom[13108] = 'b101001111;assign rom[13109] = 'b000111010;assign rom[13110] = 'b101110110;assign rom[13111] = 'b101100010;assign rom[13112] = 'b101001100;assign rom[13113] = 'b001001010;assign rom[13114] = 'b111011010;assign rom[13115] = 'b111011010;assign rom[13116] = 'b111011010;assign rom[13117] = 'b111011010;assign rom[13118] = 'b111011000;assign rom[13119] = 'b111011000;assign rom[13120] = 'b111011000;assign rom[13121] = 'b111011000;assign rom[13122] = 'b101111000;assign rom[13123] = 'b000110011;assign rom[13124] = 'b110000010;assign rom[13125] = 'b001101010;assign rom[13126] = 'b001011000;assign rom[13127] = 'b101001000;assign rom[13128] = 'b000101011;assign rom[13129] = 'b110000010;assign rom[13130] = 'b111000000;assign rom[13131] = 'b101001100;assign rom[13132] = 'b001001010;assign rom[13133] = 'b111111000;assign rom[13134] = 'b111101000;assign rom[13135] = 'b101001111;assign rom[13136] = 'b000111010;assign rom[13137] = 'b101110110;assign rom[13138] = 'b101100010;assign rom[13139] = 'b101001100;assign rom[13140] = 'b001001010;assign rom[13141] = 'b111011010;assign rom[13142] = 'b111011010;assign rom[13143] = 'b111011010;assign rom[13144] = 'b111011010;assign rom[13145] = 'b111011000;assign rom[13146] = 'b111011000;assign rom[13147] = 'b111011000;assign rom[13148] = 'b111011000;assign rom[13149] = 'b101111000;assign rom[13150] = 'b000110011;assign rom[13151] = 'b110000010;assign rom[13152] = 'b001101010;assign rom[13153] = 'b001011000;assign rom[13154] = 'b101001000;assign rom[13155] = 'b000101011;assign rom[13156] = 'b110000010;assign rom[13157] = 'b111000000;assign rom[13158] = 'b101001100;assign rom[13159] = 'b001001010;assign rom[13160] = 'b111111000;assign rom[13161] = 'b111101000;assign rom[13162] = 'b101001111;assign rom[13163] = 'b000111010;assign rom[13164] = 'b101110110;assign rom[13165] = 'b101100010;assign rom[13166] = 'b101001100;assign rom[13167] = 'b001001010;assign rom[13168] = 'b111011010;assign rom[13169] = 'b111011010;assign rom[13170] = 'b111011010;assign rom[13171] = 'b111011010;assign rom[13172] = 'b111011000;assign rom[13173] = 'b111011000;assign rom[13174] = 'b111011000;assign rom[13175] = 'b111011000;assign rom[13176] = 'b101111000;assign rom[13177] = 'b000110011;assign rom[13178] = 'b110000010;assign rom[13179] = 'b001101010;assign rom[13180] = 'b001011000;assign rom[13181] = 'b101001000;assign rom[13182] = 'b000101011;assign rom[13183] = 'b110000010;assign rom[13184] = 'b111000000;assign rom[13185] = 'b101001100;assign rom[13186] = 'b001001010;assign rom[13187] = 'b111111000;assign rom[13188] = 'b111101000;assign rom[13189] = 'b101001111;assign rom[13190] = 'b000111010;assign rom[13191] = 'b101110110;assign rom[13192] = 'b101100010;assign rom[13193] = 'b101001100;assign rom[13194] = 'b001001010;assign rom[13195] = 'b111011010;assign rom[13196] = 'b111011010;assign rom[13197] = 'b111011010;assign rom[13198] = 'b111011010;assign rom[13199] = 'b111011000;assign rom[13200] = 'b111011000;assign rom[13201] = 'b111011000;assign rom[13202] = 'b111011000;assign rom[13203] = 'b101111000;assign rom[13204] = 'b000110011;assign rom[13205] = 'b110000010;assign rom[13206] = 'b001101010;assign rom[13207] = 'b001011000;assign rom[13208] = 'b101001000;assign rom[13209] = 'b000101011;assign rom[13210] = 'b110000010;assign rom[13211] = 'b111000000;assign rom[13212] = 'b101001100;assign rom[13213] = 'b001001010;assign rom[13214] = 'b111111000;assign rom[13215] = 'b111101000;assign rom[13216] = 'b101001111;assign rom[13217] = 'b000111010;assign rom[13218] = 'b101110110;assign rom[13219] = 'b101100010;assign rom[13220] = 'b101001100;assign rom[13221] = 'b001001010;assign rom[13222] = 'b111011010;assign rom[13223] = 'b111011010;assign rom[13224] = 'b111011010;assign rom[13225] = 'b111011010;assign rom[13226] = 'b111011000;assign rom[13227] = 'b111011000;assign rom[13228] = 'b111011000;assign rom[13229] = 'b111011000;assign rom[13230] = 'b101111000;assign rom[13231] = 'b000110011;assign rom[13232] = 'b110000010;assign rom[13233] = 'b001101010;assign rom[13234] = 'b001011000;assign rom[13235] = 'b101001000;assign rom[13236] = 'b000101011;assign rom[13237] = 'b110000010;assign rom[13238] = 'b111000000;assign rom[13239] = 'b101001100;assign rom[13240] = 'b001001010;assign rom[13241] = 'b001000110;assign rom[13242] = 'b001100100;assign rom[13243] = 'b101100010;assign rom[13244] = 'b101001100;assign rom[13245] = 'b001001010;assign rom[13246] = 'b111011010;assign rom[13247] = 'b111011010;assign rom[13248] = 'b111011010;assign rom[13249] = 'b111011010;assign rom[13250] = 'b111011000;assign rom[13251] = 'b111011000;assign rom[13252] = 'b111011000;assign rom[13253] = 'b111011000;assign rom[13254] = 'b101111000;assign rom[13255] = 'b000110011;assign rom[13256] = 'b110000010;assign rom[13257] = 'b001101010;assign rom[13258] = 'b001011000;assign rom[13259] = 'b101001000;assign rom[13260] = 'b000101011;assign rom[13261] = 'b110000010;assign rom[13262] = 'b111000000;assign rom[13263] = 'b101001100;assign rom[13264] = 'b001001010;assign rom[13265] = 'b111111000;assign rom[13266] = 'b111101000;assign rom[13267] = 'b101001111;assign rom[13268] = 'b000111010;assign rom[13269] = 'b101110110;assign rom[13270] = 'b101100010;assign rom[13271] = 'b101001100;assign rom[13272] = 'b001001010;assign rom[13273] = 'b111011010;assign rom[13274] = 'b111011010;assign rom[13275] = 'b111011010;assign rom[13276] = 'b111011010;assign rom[13277] = 'b111011000;assign rom[13278] = 'b111011000;assign rom[13279] = 'b111011000;assign rom[13280] = 'b111011000;assign rom[13281] = 'b101111000;assign rom[13282] = 'b000110011;assign rom[13283] = 'b110000010;assign rom[13284] = 'b001101010;assign rom[13285] = 'b001011000;assign rom[13286] = 'b101001000;assign rom[13287] = 'b000101011;assign rom[13288] = 'b110000010;assign rom[13289] = 'b111000000;assign rom[13290] = 'b101001100;assign rom[13291] = 'b001001010;assign rom[13292] = 'b111111000;assign rom[13293] = 'b111101000;assign rom[13294] = 'b101001111;assign rom[13295] = 'b000111010;assign rom[13296] = 'b101110110;assign rom[13297] = 'b101100010;assign rom[13298] = 'b101001100;assign rom[13299] = 'b001001010;assign rom[13300] = 'b111011010;assign rom[13301] = 'b111011010;assign rom[13302] = 'b111011010;assign rom[13303] = 'b111011010;assign rom[13304] = 'b111011000;assign rom[13305] = 'b111011000;assign rom[13306] = 'b111011000;assign rom[13307] = 'b111011000;assign rom[13308] = 'b101111000;assign rom[13309] = 'b000110011;assign rom[13310] = 'b110000010;assign rom[13311] = 'b001101010;assign rom[13312] = 'b001011000;assign rom[13313] = 'b101001000;assign rom[13314] = 'b000101011;assign rom[13315] = 'b110000010;assign rom[13316] = 'b111000000;assign rom[13317] = 'b101001100;assign rom[13318] = 'b001001010;assign rom[13319] = 'b111111000;assign rom[13320] = 'b111101000;assign rom[13321] = 'b101001111;assign rom[13322] = 'b000111010;assign rom[13323] = 'b101110110;assign rom[13324] = 'b101100010;assign rom[13325] = 'b101001100;assign rom[13326] = 'b001001010;assign rom[13327] = 'b111011010;assign rom[13328] = 'b111011010;assign rom[13329] = 'b111011010;assign rom[13330] = 'b111011010;assign rom[13331] = 'b111011000;assign rom[13332] = 'b111011000;assign rom[13333] = 'b111011000;assign rom[13334] = 'b111011000;assign rom[13335] = 'b101111000;assign rom[13336] = 'b000110011;assign rom[13337] = 'b110000010;assign rom[13338] = 'b001101010;assign rom[13339] = 'b001011000;assign rom[13340] = 'b101001000;assign rom[13341] = 'b000101011;assign rom[13342] = 'b110000010;assign rom[13343] = 'b111000000;assign rom[13344] = 'b101001100;assign rom[13345] = 'b001001010;assign rom[13346] = 'b111111000;assign rom[13347] = 'b111101000;assign rom[13348] = 'b101001111;assign rom[13349] = 'b000111010;assign rom[13350] = 'b101110110;assign rom[13351] = 'b101100010;assign rom[13352] = 'b101001100;assign rom[13353] = 'b001001010;assign rom[13354] = 'b111011010;assign rom[13355] = 'b111011010;assign rom[13356] = 'b111011010;assign rom[13357] = 'b111011010;assign rom[13358] = 'b111011000;assign rom[13359] = 'b111011000;assign rom[13360] = 'b111011000;assign rom[13361] = 'b111011000;assign rom[13362] = 'b101111000;assign rom[13363] = 'b000110011;assign rom[13364] = 'b110000010;assign rom[13365] = 'b001101010;assign rom[13366] = 'b001011000;assign rom[13367] = 'b101001000;assign rom[13368] = 'b000101011;assign rom[13369] = 'b110000010;assign rom[13370] = 'b111000000;assign rom[13371] = 'b101001100;assign rom[13372] = 'b001001010;assign rom[13373] = 'b111111000;assign rom[13374] = 'b111101000;assign rom[13375] = 'b101001111;assign rom[13376] = 'b000111010;assign rom[13377] = 'b101110110;assign rom[13378] = 'b101100010;assign rom[13379] = 'b101001100;assign rom[13380] = 'b001001010;assign rom[13381] = 'b111011010;assign rom[13382] = 'b111011010;assign rom[13383] = 'b111011010;assign rom[13384] = 'b111011010;assign rom[13385] = 'b111011000;assign rom[13386] = 'b111011000;assign rom[13387] = 'b111011000;assign rom[13388] = 'b111011000;assign rom[13389] = 'b101111000;assign rom[13390] = 'b000110011;assign rom[13391] = 'b110000010;assign rom[13392] = 'b001101010;assign rom[13393] = 'b001011000;assign rom[13394] = 'b101001000;assign rom[13395] = 'b000101011;assign rom[13396] = 'b110000010;assign rom[13397] = 'b111000000;assign rom[13398] = 'b101001100;assign rom[13399] = 'b001001010;assign rom[13400] = 'b111111000;assign rom[13401] = 'b111101000;assign rom[13402] = 'b101001111;assign rom[13403] = 'b000111010;assign rom[13404] = 'b101110110;assign rom[13405] = 'b101100010;assign rom[13406] = 'b101001100;assign rom[13407] = 'b001001010;assign rom[13408] = 'b111011010;assign rom[13409] = 'b111011010;assign rom[13410] = 'b111011010;assign rom[13411] = 'b111011010;assign rom[13412] = 'b111011000;assign rom[13413] = 'b111011000;assign rom[13414] = 'b111011000;assign rom[13415] = 'b111011000;assign rom[13416] = 'b101111000;assign rom[13417] = 'b000110011;assign rom[13418] = 'b110000010;assign rom[13419] = 'b001101010;assign rom[13420] = 'b001011000;assign rom[13421] = 'b101001000;assign rom[13422] = 'b000101011;assign rom[13423] = 'b110000010;assign rom[13424] = 'b111000000;assign rom[13425] = 'b101001100;assign rom[13426] = 'b001001010;assign rom[13427] = 'b111111000;assign rom[13428] = 'b111101000;assign rom[13429] = 'b101001111;assign rom[13430] = 'b000111010;assign rom[13431] = 'b101110110;assign rom[13432] = 'b101100010;assign rom[13433] = 'b101001100;assign rom[13434] = 'b001001010;assign rom[13435] = 'b111011010;assign rom[13436] = 'b111011010;assign rom[13437] = 'b111011010;assign rom[13438] = 'b111011010;assign rom[13439] = 'b111011000;assign rom[13440] = 'b111011000;assign rom[13441] = 'b111011000;assign rom[13442] = 'b111011000;assign rom[13443] = 'b101111000;assign rom[13444] = 'b000110011;assign rom[13445] = 'b110000010;assign rom[13446] = 'b001101010;assign rom[13447] = 'b001011000;assign rom[13448] = 'b101001000;assign rom[13449] = 'b000101011;assign rom[13450] = 'b110000010;assign rom[13451] = 'b111000000;assign rom[13452] = 'b101001100;assign rom[13453] = 'b001001010;assign rom[13454] = 'b111111000;assign rom[13455] = 'b111101000;assign rom[13456] = 'b101001111;assign rom[13457] = 'b000111010;assign rom[13458] = 'b101110110;assign rom[13459] = 'b101100010;assign rom[13460] = 'b101001100;assign rom[13461] = 'b001001010;assign rom[13462] = 'b111011010;assign rom[13463] = 'b111011010;assign rom[13464] = 'b111011010;assign rom[13465] = 'b111011010;assign rom[13466] = 'b111011000;assign rom[13467] = 'b111011000;assign rom[13468] = 'b111011000;assign rom[13469] = 'b111011000;assign rom[13470] = 'b101111000;assign rom[13471] = 'b000110011;assign rom[13472] = 'b110000010;assign rom[13473] = 'b001101010;assign rom[13474] = 'b001011000;assign rom[13475] = 'b101001000;assign rom[13476] = 'b000101011;assign rom[13477] = 'b110000010;assign rom[13478] = 'b111000000;assign rom[13479] = 'b101001100;assign rom[13480] = 'b001001010;assign rom[13481] = 'b001000110;assign rom[13482] = 'b001100100;assign rom[13483] = 'b101100010;assign rom[13484] = 'b101001100;assign rom[13485] = 'b001001010;assign rom[13486] = 'b111011010;assign rom[13487] = 'b111011010;assign rom[13488] = 'b111011010;assign rom[13489] = 'b111011010;assign rom[13490] = 'b111011000;assign rom[13491] = 'b111011000;assign rom[13492] = 'b111011000;assign rom[13493] = 'b111011000;assign rom[13494] = 'b101111000;assign rom[13495] = 'b000110011;assign rom[13496] = 'b110000010;assign rom[13497] = 'b001101010;assign rom[13498] = 'b001011000;assign rom[13499] = 'b101001000;assign rom[13500] = 'b000101011;assign rom[13501] = 'b110000010;assign rom[13502] = 'b111000000;assign rom[13503] = 'b101001100;assign rom[13504] = 'b001001010;assign rom[13505] = 'b111111000;assign rom[13506] = 'b111101000;assign rom[13507] = 'b101001111;assign rom[13508] = 'b000111010;assign rom[13509] = 'b101110110;assign rom[13510] = 'b101100010;assign rom[13511] = 'b101001100;assign rom[13512] = 'b001001010;assign rom[13513] = 'b111011010;assign rom[13514] = 'b111011010;assign rom[13515] = 'b111011010;assign rom[13516] = 'b111011010;assign rom[13517] = 'b111011000;assign rom[13518] = 'b111011000;assign rom[13519] = 'b111011000;assign rom[13520] = 'b111011000;assign rom[13521] = 'b101111000;assign rom[13522] = 'b000110011;assign rom[13523] = 'b110000010;assign rom[13524] = 'b001101010;assign rom[13525] = 'b001011000;assign rom[13526] = 'b101001000;assign rom[13527] = 'b000101011;assign rom[13528] = 'b110000010;assign rom[13529] = 'b111000000;assign rom[13530] = 'b101001100;assign rom[13531] = 'b001001010;assign rom[13532] = 'b111111000;assign rom[13533] = 'b111101000;assign rom[13534] = 'b101001111;assign rom[13535] = 'b000111010;assign rom[13536] = 'b101110110;assign rom[13537] = 'b101100010;assign rom[13538] = 'b101001100;assign rom[13539] = 'b001001010;assign rom[13540] = 'b111011010;assign rom[13541] = 'b111011010;assign rom[13542] = 'b111011010;assign rom[13543] = 'b111011010;assign rom[13544] = 'b111011000;assign rom[13545] = 'b111011000;assign rom[13546] = 'b111011000;assign rom[13547] = 'b111011000;assign rom[13548] = 'b101111000;assign rom[13549] = 'b000110011;assign rom[13550] = 'b110000010;assign rom[13551] = 'b001101010;assign rom[13552] = 'b001011000;assign rom[13553] = 'b101001000;assign rom[13554] = 'b000101011;assign rom[13555] = 'b110000010;assign rom[13556] = 'b111000000;assign rom[13557] = 'b101001100;assign rom[13558] = 'b001001010;assign rom[13559] = 'b111111000;assign rom[13560] = 'b111101000;assign rom[13561] = 'b101001111;assign rom[13562] = 'b000111010;assign rom[13563] = 'b101110110;assign rom[13564] = 'b101100010;assign rom[13565] = 'b101001100;assign rom[13566] = 'b001001010;assign rom[13567] = 'b111011010;assign rom[13568] = 'b111011010;assign rom[13569] = 'b111011010;assign rom[13570] = 'b111011010;assign rom[13571] = 'b111011000;assign rom[13572] = 'b111011000;assign rom[13573] = 'b111011000;assign rom[13574] = 'b111011000;assign rom[13575] = 'b101111000;assign rom[13576] = 'b000110011;assign rom[13577] = 'b110000010;assign rom[13578] = 'b001101010;assign rom[13579] = 'b001011000;assign rom[13580] = 'b101001000;assign rom[13581] = 'b000101011;assign rom[13582] = 'b110000010;assign rom[13583] = 'b111000000;assign rom[13584] = 'b101001100;assign rom[13585] = 'b001001010;assign rom[13586] = 'b111111000;assign rom[13587] = 'b111101000;assign rom[13588] = 'b101001111;assign rom[13589] = 'b000111010;assign rom[13590] = 'b101110110;assign rom[13591] = 'b101100010;assign rom[13592] = 'b101001100;assign rom[13593] = 'b001001010;assign rom[13594] = 'b111011010;assign rom[13595] = 'b111011010;assign rom[13596] = 'b111011010;assign rom[13597] = 'b111011010;assign rom[13598] = 'b111011000;assign rom[13599] = 'b111011000;assign rom[13600] = 'b111011000;assign rom[13601] = 'b111011000;assign rom[13602] = 'b101111000;assign rom[13603] = 'b000110011;assign rom[13604] = 'b110000010;assign rom[13605] = 'b001101010;assign rom[13606] = 'b001011000;assign rom[13607] = 'b101001000;assign rom[13608] = 'b000101011;assign rom[13609] = 'b110000010;assign rom[13610] = 'b111000000;assign rom[13611] = 'b101001100;assign rom[13612] = 'b001001010;assign rom[13613] = 'b111111000;assign rom[13614] = 'b111101000;assign rom[13615] = 'b101001111;assign rom[13616] = 'b000111010;assign rom[13617] = 'b101110110;assign rom[13618] = 'b101100010;assign rom[13619] = 'b101001100;assign rom[13620] = 'b001001010;assign rom[13621] = 'b111011010;assign rom[13622] = 'b111011010;assign rom[13623] = 'b111011010;assign rom[13624] = 'b111011010;assign rom[13625] = 'b111011000;assign rom[13626] = 'b111011000;assign rom[13627] = 'b111011000;assign rom[13628] = 'b111011000;assign rom[13629] = 'b101111000;assign rom[13630] = 'b000110011;assign rom[13631] = 'b110000010;assign rom[13632] = 'b001101010;assign rom[13633] = 'b001011000;assign rom[13634] = 'b101001000;assign rom[13635] = 'b000101011;assign rom[13636] = 'b110000010;assign rom[13637] = 'b111000000;assign rom[13638] = 'b101001100;assign rom[13639] = 'b001001010;assign rom[13640] = 'b111111000;assign rom[13641] = 'b111101000;assign rom[13642] = 'b101001111;assign rom[13643] = 'b000111010;assign rom[13644] = 'b101110110;assign rom[13645] = 'b101100010;assign rom[13646] = 'b101001100;assign rom[13647] = 'b001001010;assign rom[13648] = 'b111011010;assign rom[13649] = 'b111011010;assign rom[13650] = 'b111011010;assign rom[13651] = 'b111011010;assign rom[13652] = 'b111011000;assign rom[13653] = 'b111011000;assign rom[13654] = 'b111011000;assign rom[13655] = 'b111011000;assign rom[13656] = 'b101111000;assign rom[13657] = 'b000110011;assign rom[13658] = 'b110000010;assign rom[13659] = 'b001101010;assign rom[13660] = 'b001011000;assign rom[13661] = 'b101001000;assign rom[13662] = 'b000101011;assign rom[13663] = 'b110000010;assign rom[13664] = 'b111000000;assign rom[13665] = 'b101001100;assign rom[13666] = 'b001001010;assign rom[13667] = 'b111111000;assign rom[13668] = 'b111101000;assign rom[13669] = 'b101001111;assign rom[13670] = 'b000111010;assign rom[13671] = 'b101110110;assign rom[13672] = 'b101100010;assign rom[13673] = 'b101001100;assign rom[13674] = 'b001001010;assign rom[13675] = 'b111011010;assign rom[13676] = 'b111011010;assign rom[13677] = 'b111011010;assign rom[13678] = 'b111011010;assign rom[13679] = 'b111011000;assign rom[13680] = 'b111011000;assign rom[13681] = 'b111011000;assign rom[13682] = 'b111011000;assign rom[13683] = 'b101111000;assign rom[13684] = 'b000110011;assign rom[13685] = 'b110000010;assign rom[13686] = 'b001101010;assign rom[13687] = 'b001011000;assign rom[13688] = 'b101001000;assign rom[13689] = 'b000101011;assign rom[13690] = 'b110000010;assign rom[13691] = 'b111000000;assign rom[13692] = 'b101001100;assign rom[13693] = 'b001001010;assign rom[13694] = 'b111111000;assign rom[13695] = 'b111101000;assign rom[13696] = 'b101001111;assign rom[13697] = 'b000111010;assign rom[13698] = 'b101110110;assign rom[13699] = 'b101100010;assign rom[13700] = 'b101001100;assign rom[13701] = 'b001001010;assign rom[13702] = 'b111011010;assign rom[13703] = 'b111011010;assign rom[13704] = 'b111011010;assign rom[13705] = 'b111011010;assign rom[13706] = 'b111011000;assign rom[13707] = 'b111011000;assign rom[13708] = 'b111011000;assign rom[13709] = 'b111011000;assign rom[13710] = 'b101111000;assign rom[13711] = 'b000110011;assign rom[13712] = 'b110000010;assign rom[13713] = 'b001101010;assign rom[13714] = 'b001011000;assign rom[13715] = 'b101001000;assign rom[13716] = 'b000101011;assign rom[13717] = 'b110000010;assign rom[13718] = 'b111000000;assign rom[13719] = 'b101001100;assign rom[13720] = 'b001001010;assign rom[13721] = 'b001000110;assign rom[13722] = 'b001100100;assign rom[13723] = 'b101100010;assign rom[13724] = 'b101001100;assign rom[13725] = 'b001001010;assign rom[13726] = 'b111011010;assign rom[13727] = 'b111011010;assign rom[13728] = 'b111011010;assign rom[13729] = 'b111011010;assign rom[13730] = 'b111011000;assign rom[13731] = 'b111011000;assign rom[13732] = 'b111011000;assign rom[13733] = 'b111011000;assign rom[13734] = 'b101111000;assign rom[13735] = 'b000110011;assign rom[13736] = 'b110000010;assign rom[13737] = 'b001101010;assign rom[13738] = 'b001011000;assign rom[13739] = 'b101001000;assign rom[13740] = 'b000101011;assign rom[13741] = 'b110000010;assign rom[13742] = 'b111000000;assign rom[13743] = 'b101001100;assign rom[13744] = 'b001001010;assign rom[13745] = 'b111111000;assign rom[13746] = 'b111101000;assign rom[13747] = 'b101001111;assign rom[13748] = 'b000111010;assign rom[13749] = 'b101110110;assign rom[13750] = 'b101100010;assign rom[13751] = 'b101001100;assign rom[13752] = 'b001001010;assign rom[13753] = 'b111011010;assign rom[13754] = 'b111011010;assign rom[13755] = 'b111011010;assign rom[13756] = 'b111011010;assign rom[13757] = 'b111011000;assign rom[13758] = 'b111011000;assign rom[13759] = 'b111011000;assign rom[13760] = 'b111011000;assign rom[13761] = 'b101111000;assign rom[13762] = 'b000110011;assign rom[13763] = 'b110000010;assign rom[13764] = 'b001101010;assign rom[13765] = 'b001011000;assign rom[13766] = 'b101001000;assign rom[13767] = 'b000101011;assign rom[13768] = 'b110000010;assign rom[13769] = 'b111000000;assign rom[13770] = 'b101001100;assign rom[13771] = 'b001001010;assign rom[13772] = 'b111111000;assign rom[13773] = 'b111101000;assign rom[13774] = 'b101001111;assign rom[13775] = 'b000111010;assign rom[13776] = 'b101110110;assign rom[13777] = 'b101100010;assign rom[13778] = 'b101001100;assign rom[13779] = 'b001001010;assign rom[13780] = 'b111011010;assign rom[13781] = 'b111011010;assign rom[13782] = 'b111011010;assign rom[13783] = 'b111011010;assign rom[13784] = 'b111011000;assign rom[13785] = 'b111011000;assign rom[13786] = 'b111011000;assign rom[13787] = 'b111011000;assign rom[13788] = 'b101111000;assign rom[13789] = 'b000110011;assign rom[13790] = 'b110000010;assign rom[13791] = 'b001101010;assign rom[13792] = 'b001011000;assign rom[13793] = 'b101001000;assign rom[13794] = 'b000101011;assign rom[13795] = 'b110000010;assign rom[13796] = 'b111000000;assign rom[13797] = 'b101001100;assign rom[13798] = 'b001001010;assign rom[13799] = 'b111111000;assign rom[13800] = 'b111101000;assign rom[13801] = 'b101001111;assign rom[13802] = 'b000111010;assign rom[13803] = 'b101110110;assign rom[13804] = 'b101100010;assign rom[13805] = 'b101001100;assign rom[13806] = 'b001001010;assign rom[13807] = 'b111011010;assign rom[13808] = 'b111011010;assign rom[13809] = 'b111011010;assign rom[13810] = 'b111011010;assign rom[13811] = 'b111011000;assign rom[13812] = 'b111011000;assign rom[13813] = 'b111011000;assign rom[13814] = 'b111011000;assign rom[13815] = 'b101111000;assign rom[13816] = 'b000110011;assign rom[13817] = 'b110000010;assign rom[13818] = 'b001101010;assign rom[13819] = 'b001011000;assign rom[13820] = 'b101001000;assign rom[13821] = 'b000101011;assign rom[13822] = 'b110000010;assign rom[13823] = 'b111000000;assign rom[13824] = 'b101001100;assign rom[13825] = 'b001001010;assign rom[13826] = 'b111111000;assign rom[13827] = 'b111101000;assign rom[13828] = 'b101001111;assign rom[13829] = 'b000111010;assign rom[13830] = 'b101110110;assign rom[13831] = 'b101100010;assign rom[13832] = 'b101001100;assign rom[13833] = 'b001001010;assign rom[13834] = 'b111011010;assign rom[13835] = 'b111011010;assign rom[13836] = 'b111011010;assign rom[13837] = 'b111011010;assign rom[13838] = 'b111011000;assign rom[13839] = 'b111011000;assign rom[13840] = 'b111011000;assign rom[13841] = 'b111011000;assign rom[13842] = 'b101111000;assign rom[13843] = 'b000110011;assign rom[13844] = 'b110000010;assign rom[13845] = 'b001101010;assign rom[13846] = 'b001011000;assign rom[13847] = 'b101001000;assign rom[13848] = 'b000101011;assign rom[13849] = 'b110000010;assign rom[13850] = 'b111000000;assign rom[13851] = 'b101001100;assign rom[13852] = 'b001001010;assign rom[13853] = 'b111111000;assign rom[13854] = 'b111101000;assign rom[13855] = 'b101001111;assign rom[13856] = 'b000111010;assign rom[13857] = 'b101110110;assign rom[13858] = 'b101100010;assign rom[13859] = 'b101001100;assign rom[13860] = 'b001001010;assign rom[13861] = 'b111011010;assign rom[13862] = 'b111011010;assign rom[13863] = 'b111011010;assign rom[13864] = 'b111011010;assign rom[13865] = 'b111011000;assign rom[13866] = 'b111011000;assign rom[13867] = 'b111011000;assign rom[13868] = 'b111011000;assign rom[13869] = 'b101111000;assign rom[13870] = 'b000110011;assign rom[13871] = 'b110000010;assign rom[13872] = 'b001101010;assign rom[13873] = 'b001011000;assign rom[13874] = 'b101001000;assign rom[13875] = 'b000101011;assign rom[13876] = 'b110000010;assign rom[13877] = 'b111000000;assign rom[13878] = 'b101001100;assign rom[13879] = 'b001001010;assign rom[13880] = 'b111111000;assign rom[13881] = 'b111101000;assign rom[13882] = 'b101001111;assign rom[13883] = 'b000111010;assign rom[13884] = 'b101110110;assign rom[13885] = 'b101100010;assign rom[13886] = 'b101001100;assign rom[13887] = 'b001001010;assign rom[13888] = 'b111011010;assign rom[13889] = 'b111011010;assign rom[13890] = 'b111011010;assign rom[13891] = 'b111011010;assign rom[13892] = 'b111011000;assign rom[13893] = 'b111011000;assign rom[13894] = 'b111011000;assign rom[13895] = 'b111011000;assign rom[13896] = 'b101111000;assign rom[13897] = 'b000110011;assign rom[13898] = 'b110000010;assign rom[13899] = 'b001101010;assign rom[13900] = 'b001011000;assign rom[13901] = 'b101001000;assign rom[13902] = 'b000101011;assign rom[13903] = 'b110000010;assign rom[13904] = 'b111000000;assign rom[13905] = 'b101001100;assign rom[13906] = 'b001001010;assign rom[13907] = 'b111111000;assign rom[13908] = 'b111101000;assign rom[13909] = 'b101001111;assign rom[13910] = 'b000111010;assign rom[13911] = 'b101110110;assign rom[13912] = 'b101100010;assign rom[13913] = 'b101001100;assign rom[13914] = 'b001001010;assign rom[13915] = 'b111011010;assign rom[13916] = 'b111011010;assign rom[13917] = 'b111011010;assign rom[13918] = 'b111011010;assign rom[13919] = 'b111011000;assign rom[13920] = 'b111011000;assign rom[13921] = 'b111011000;assign rom[13922] = 'b111011000;assign rom[13923] = 'b101111000;assign rom[13924] = 'b000110011;assign rom[13925] = 'b110000010;assign rom[13926] = 'b001101010;assign rom[13927] = 'b001011000;assign rom[13928] = 'b101001000;assign rom[13929] = 'b000101011;assign rom[13930] = 'b110000010;assign rom[13931] = 'b111000000;assign rom[13932] = 'b101001100;assign rom[13933] = 'b001001010;assign rom[13934] = 'b111111000;assign rom[13935] = 'b111101000;assign rom[13936] = 'b101001111;assign rom[13937] = 'b000111010;assign rom[13938] = 'b101110110;assign rom[13939] = 'b101100010;assign rom[13940] = 'b101001100;assign rom[13941] = 'b001001010;assign rom[13942] = 'b111011010;assign rom[13943] = 'b111011010;assign rom[13944] = 'b111011010;assign rom[13945] = 'b111011010;assign rom[13946] = 'b111011000;assign rom[13947] = 'b111011000;assign rom[13948] = 'b111011000;assign rom[13949] = 'b111011000;assign rom[13950] = 'b101111000;assign rom[13951] = 'b000110011;assign rom[13952] = 'b110000010;assign rom[13953] = 'b001101010;assign rom[13954] = 'b001011000;assign rom[13955] = 'b101001000;assign rom[13956] = 'b000101011;assign rom[13957] = 'b110000010;assign rom[13958] = 'b111000000;assign rom[13959] = 'b101001100;assign rom[13960] = 'b001001010;assign rom[13961] = 'b001000110;assign rom[13962] = 'b001100100;assign rom[13963] = 'b101100010;assign rom[13964] = 'b101001100;assign rom[13965] = 'b001001010;assign rom[13966] = 'b111011010;assign rom[13967] = 'b111011010;assign rom[13968] = 'b111011010;assign rom[13969] = 'b111011010;assign rom[13970] = 'b111011000;assign rom[13971] = 'b111011000;assign rom[13972] = 'b111011000;assign rom[13973] = 'b111011000;assign rom[13974] = 'b101111000;assign rom[13975] = 'b000110011;assign rom[13976] = 'b110000010;assign rom[13977] = 'b001101010;assign rom[13978] = 'b001011000;assign rom[13979] = 'b101001000;assign rom[13980] = 'b000101011;assign rom[13981] = 'b110000010;assign rom[13982] = 'b111000000;assign rom[13983] = 'b101001100;assign rom[13984] = 'b001001010;assign rom[13985] = 'b111111000;assign rom[13986] = 'b111101000;assign rom[13987] = 'b101001111;assign rom[13988] = 'b000111010;assign rom[13989] = 'b101110110;assign rom[13990] = 'b101100010;assign rom[13991] = 'b101001100;assign rom[13992] = 'b001001010;assign rom[13993] = 'b111011010;assign rom[13994] = 'b111011010;assign rom[13995] = 'b111011010;assign rom[13996] = 'b111011010;assign rom[13997] = 'b111011000;assign rom[13998] = 'b111011000;assign rom[13999] = 'b111011000;assign rom[14000] = 'b111011000;assign rom[14001] = 'b101111000;assign rom[14002] = 'b000110011;assign rom[14003] = 'b110000010;assign rom[14004] = 'b001101010;assign rom[14005] = 'b001011000;assign rom[14006] = 'b101001000;assign rom[14007] = 'b000101011;assign rom[14008] = 'b110000010;assign rom[14009] = 'b111000000;assign rom[14010] = 'b101001100;assign rom[14011] = 'b001001010;assign rom[14012] = 'b111111000;assign rom[14013] = 'b111101000;assign rom[14014] = 'b101001111;assign rom[14015] = 'b000111010;assign rom[14016] = 'b101110110;assign rom[14017] = 'b101100010;assign rom[14018] = 'b101001100;assign rom[14019] = 'b001001010;assign rom[14020] = 'b111011010;assign rom[14021] = 'b111011010;assign rom[14022] = 'b111011010;assign rom[14023] = 'b111011010;assign rom[14024] = 'b111011000;assign rom[14025] = 'b111011000;assign rom[14026] = 'b111011000;assign rom[14027] = 'b111011000;assign rom[14028] = 'b101111000;assign rom[14029] = 'b000110011;assign rom[14030] = 'b110000010;assign rom[14031] = 'b001101010;assign rom[14032] = 'b001011000;assign rom[14033] = 'b101001000;assign rom[14034] = 'b000101011;assign rom[14035] = 'b110000010;assign rom[14036] = 'b111000000;assign rom[14037] = 'b101001100;assign rom[14038] = 'b001001010;assign rom[14039] = 'b111111000;assign rom[14040] = 'b111101000;assign rom[14041] = 'b101001111;assign rom[14042] = 'b000111010;assign rom[14043] = 'b101110110;assign rom[14044] = 'b101100010;assign rom[14045] = 'b101001100;assign rom[14046] = 'b001001010;assign rom[14047] = 'b111011010;assign rom[14048] = 'b111011010;assign rom[14049] = 'b111011010;assign rom[14050] = 'b111011010;assign rom[14051] = 'b111011000;assign rom[14052] = 'b111011000;assign rom[14053] = 'b111011000;assign rom[14054] = 'b111011000;assign rom[14055] = 'b101111000;assign rom[14056] = 'b000110011;assign rom[14057] = 'b110000010;assign rom[14058] = 'b001101010;assign rom[14059] = 'b001011000;assign rom[14060] = 'b101001000;assign rom[14061] = 'b000101011;assign rom[14062] = 'b110000010;assign rom[14063] = 'b111000000;assign rom[14064] = 'b101001100;assign rom[14065] = 'b001001010;assign rom[14066] = 'b111111000;assign rom[14067] = 'b111101000;assign rom[14068] = 'b101001111;assign rom[14069] = 'b000111010;assign rom[14070] = 'b101110110;assign rom[14071] = 'b101100010;assign rom[14072] = 'b101001100;assign rom[14073] = 'b001001010;assign rom[14074] = 'b111011010;assign rom[14075] = 'b111011010;assign rom[14076] = 'b111011010;assign rom[14077] = 'b111011010;assign rom[14078] = 'b111011000;assign rom[14079] = 'b111011000;assign rom[14080] = 'b111011000;assign rom[14081] = 'b111011000;assign rom[14082] = 'b101111000;assign rom[14083] = 'b000110011;assign rom[14084] = 'b110000010;assign rom[14085] = 'b001101010;assign rom[14086] = 'b001011000;assign rom[14087] = 'b101001000;assign rom[14088] = 'b000101011;assign rom[14089] = 'b110000010;assign rom[14090] = 'b111000000;assign rom[14091] = 'b101001100;assign rom[14092] = 'b001001010;assign rom[14093] = 'b111111000;assign rom[14094] = 'b111101000;assign rom[14095] = 'b101001111;assign rom[14096] = 'b000111010;assign rom[14097] = 'b101110110;assign rom[14098] = 'b101100010;assign rom[14099] = 'b101001100;assign rom[14100] = 'b001001010;assign rom[14101] = 'b111011010;assign rom[14102] = 'b111011010;assign rom[14103] = 'b111011010;assign rom[14104] = 'b111011010;assign rom[14105] = 'b111011000;assign rom[14106] = 'b111011000;assign rom[14107] = 'b111011000;assign rom[14108] = 'b111011000;assign rom[14109] = 'b101111000;assign rom[14110] = 'b000110011;assign rom[14111] = 'b110000010;assign rom[14112] = 'b001101010;assign rom[14113] = 'b001011000;assign rom[14114] = 'b101001000;assign rom[14115] = 'b000101011;assign rom[14116] = 'b110000010;assign rom[14117] = 'b111000000;assign rom[14118] = 'b101001100;assign rom[14119] = 'b001001010;assign rom[14120] = 'b111111000;assign rom[14121] = 'b111101000;assign rom[14122] = 'b101001111;assign rom[14123] = 'b000111010;assign rom[14124] = 'b101110110;assign rom[14125] = 'b101100010;assign rom[14126] = 'b101001100;assign rom[14127] = 'b001001010;assign rom[14128] = 'b111011010;assign rom[14129] = 'b111011010;assign rom[14130] = 'b111011010;assign rom[14131] = 'b111011010;assign rom[14132] = 'b111011000;assign rom[14133] = 'b111011000;assign rom[14134] = 'b111011000;assign rom[14135] = 'b111011000;assign rom[14136] = 'b101111000;assign rom[14137] = 'b000110011;assign rom[14138] = 'b110000010;assign rom[14139] = 'b001101010;assign rom[14140] = 'b001011000;assign rom[14141] = 'b101001000;assign rom[14142] = 'b000101011;assign rom[14143] = 'b110000010;assign rom[14144] = 'b111000000;assign rom[14145] = 'b101001100;assign rom[14146] = 'b001001010;assign rom[14147] = 'b111111000;assign rom[14148] = 'b111101000;assign rom[14149] = 'b101001111;assign rom[14150] = 'b000111010;assign rom[14151] = 'b101110110;assign rom[14152] = 'b101100010;assign rom[14153] = 'b101001100;assign rom[14154] = 'b001001010;assign rom[14155] = 'b111011010;assign rom[14156] = 'b111011010;assign rom[14157] = 'b111011010;assign rom[14158] = 'b111011010;assign rom[14159] = 'b111011000;assign rom[14160] = 'b111011000;assign rom[14161] = 'b111011000;assign rom[14162] = 'b111011000;assign rom[14163] = 'b101111000;assign rom[14164] = 'b000110011;assign rom[14165] = 'b110000010;assign rom[14166] = 'b001101010;assign rom[14167] = 'b001011000;assign rom[14168] = 'b101001000;assign rom[14169] = 'b000101011;assign rom[14170] = 'b110000010;assign rom[14171] = 'b111000000;assign rom[14172] = 'b101001100;assign rom[14173] = 'b001001010;assign rom[14174] = 'b111111000;assign rom[14175] = 'b111101000;assign rom[14176] = 'b101001111;assign rom[14177] = 'b000111010;assign rom[14178] = 'b101110110;assign rom[14179] = 'b101100010;assign rom[14180] = 'b101001100;assign rom[14181] = 'b001001010;assign rom[14182] = 'b111011010;assign rom[14183] = 'b111011010;assign rom[14184] = 'b111011010;assign rom[14185] = 'b111011010;assign rom[14186] = 'b111011000;assign rom[14187] = 'b111011000;assign rom[14188] = 'b111011000;assign rom[14189] = 'b111011000;assign rom[14190] = 'b101111000;assign rom[14191] = 'b000110011;assign rom[14192] = 'b110000010;assign rom[14193] = 'b001101010;assign rom[14194] = 'b001011000;assign rom[14195] = 'b101001000;assign rom[14196] = 'b000101011;assign rom[14197] = 'b110000010;assign rom[14198] = 'b111000000;assign rom[14199] = 'b101001100;assign rom[14200] = 'b001001010;assign rom[14201] = 'b001000110;assign rom[14202] = 'b001100100;assign rom[14203] = 'b101100010;assign rom[14204] = 'b101001100;assign rom[14205] = 'b001001010;assign rom[14206] = 'b111011010;assign rom[14207] = 'b111011010;assign rom[14208] = 'b111011010;assign rom[14209] = 'b111011010;assign rom[14210] = 'b111011000;assign rom[14211] = 'b111011000;assign rom[14212] = 'b111011000;assign rom[14213] = 'b111011000;assign rom[14214] = 'b101111000;assign rom[14215] = 'b000110011;assign rom[14216] = 'b110000010;assign rom[14217] = 'b001101010;assign rom[14218] = 'b001011000;assign rom[14219] = 'b101001000;assign rom[14220] = 'b000101011;assign rom[14221] = 'b110000010;assign rom[14222] = 'b111000000;assign rom[14223] = 'b101001100;assign rom[14224] = 'b001001010;assign rom[14225] = 'b111111000;assign rom[14226] = 'b111101000;assign rom[14227] = 'b101001111;assign rom[14228] = 'b000111010;assign rom[14229] = 'b101110110;assign rom[14230] = 'b101100010;assign rom[14231] = 'b101001100;assign rom[14232] = 'b001001010;assign rom[14233] = 'b111011010;assign rom[14234] = 'b111011010;assign rom[14235] = 'b111011010;assign rom[14236] = 'b111011010;assign rom[14237] = 'b111011000;assign rom[14238] = 'b111011000;assign rom[14239] = 'b111011000;assign rom[14240] = 'b111011000;assign rom[14241] = 'b101111000;assign rom[14242] = 'b000110011;assign rom[14243] = 'b110000010;assign rom[14244] = 'b001101010;assign rom[14245] = 'b001011000;assign rom[14246] = 'b101001000;assign rom[14247] = 'b000101011;assign rom[14248] = 'b110000010;assign rom[14249] = 'b111000000;assign rom[14250] = 'b101001100;assign rom[14251] = 'b001001010;assign rom[14252] = 'b111111000;assign rom[14253] = 'b111101000;assign rom[14254] = 'b101001111;assign rom[14255] = 'b000111010;assign rom[14256] = 'b101110110;assign rom[14257] = 'b101100010;assign rom[14258] = 'b101001100;assign rom[14259] = 'b001001010;assign rom[14260] = 'b111011010;assign rom[14261] = 'b111011010;assign rom[14262] = 'b111011010;assign rom[14263] = 'b111011010;assign rom[14264] = 'b111011000;assign rom[14265] = 'b111011000;assign rom[14266] = 'b111011000;assign rom[14267] = 'b111011000;assign rom[14268] = 'b101111000;assign rom[14269] = 'b000110011;assign rom[14270] = 'b110000010;assign rom[14271] = 'b001101010;assign rom[14272] = 'b001011000;assign rom[14273] = 'b101001000;assign rom[14274] = 'b000101011;assign rom[14275] = 'b110000010;assign rom[14276] = 'b111000000;assign rom[14277] = 'b101001100;assign rom[14278] = 'b001001010;assign rom[14279] = 'b111111000;assign rom[14280] = 'b111101000;assign rom[14281] = 'b101001111;assign rom[14282] = 'b000111010;assign rom[14283] = 'b101110110;assign rom[14284] = 'b101100010;assign rom[14285] = 'b101001100;assign rom[14286] = 'b001001010;assign rom[14287] = 'b111011010;assign rom[14288] = 'b111011010;assign rom[14289] = 'b111011010;assign rom[14290] = 'b111011010;assign rom[14291] = 'b111011000;assign rom[14292] = 'b111011000;assign rom[14293] = 'b111011000;assign rom[14294] = 'b111011000;assign rom[14295] = 'b101111000;assign rom[14296] = 'b000110011;assign rom[14297] = 'b110000010;assign rom[14298] = 'b001101010;assign rom[14299] = 'b001011000;assign rom[14300] = 'b101001000;assign rom[14301] = 'b000101011;assign rom[14302] = 'b110000010;assign rom[14303] = 'b111000000;assign rom[14304] = 'b101001100;assign rom[14305] = 'b001001010;assign rom[14306] = 'b111111000;assign rom[14307] = 'b111101000;assign rom[14308] = 'b101001111;assign rom[14309] = 'b000111010;assign rom[14310] = 'b101110110;assign rom[14311] = 'b101100010;assign rom[14312] = 'b101001100;assign rom[14313] = 'b001001010;assign rom[14314] = 'b111011010;assign rom[14315] = 'b111011010;assign rom[14316] = 'b111011010;assign rom[14317] = 'b111011010;assign rom[14318] = 'b111011000;assign rom[14319] = 'b111011000;assign rom[14320] = 'b111011000;assign rom[14321] = 'b111011000;assign rom[14322] = 'b101111000;assign rom[14323] = 'b000110011;assign rom[14324] = 'b110000010;assign rom[14325] = 'b001101010;assign rom[14326] = 'b001011000;assign rom[14327] = 'b101001000;assign rom[14328] = 'b000101011;assign rom[14329] = 'b110000010;assign rom[14330] = 'b111000000;assign rom[14331] = 'b101001100;assign rom[14332] = 'b001001010;assign rom[14333] = 'b111111000;assign rom[14334] = 'b111101000;assign rom[14335] = 'b101001111;assign rom[14336] = 'b000111010;assign rom[14337] = 'b101110110;assign rom[14338] = 'b101100010;assign rom[14339] = 'b101001100;assign rom[14340] = 'b001001010;assign rom[14341] = 'b111011010;assign rom[14342] = 'b111011010;assign rom[14343] = 'b111011010;assign rom[14344] = 'b111011010;assign rom[14345] = 'b111011000;assign rom[14346] = 'b111011000;assign rom[14347] = 'b111011000;assign rom[14348] = 'b111011000;assign rom[14349] = 'b101111000;assign rom[14350] = 'b000110011;assign rom[14351] = 'b110000010;assign rom[14352] = 'b001101010;assign rom[14353] = 'b001011000;assign rom[14354] = 'b101001000;assign rom[14355] = 'b000101011;assign rom[14356] = 'b110000010;assign rom[14357] = 'b111000000;assign rom[14358] = 'b101001100;assign rom[14359] = 'b001001010;assign rom[14360] = 'b111111000;assign rom[14361] = 'b111101000;assign rom[14362] = 'b101001111;assign rom[14363] = 'b000111010;assign rom[14364] = 'b101110110;assign rom[14365] = 'b101100010;assign rom[14366] = 'b101001100;assign rom[14367] = 'b001001010;assign rom[14368] = 'b111011010;assign rom[14369] = 'b111011010;assign rom[14370] = 'b111011010;assign rom[14371] = 'b111011010;assign rom[14372] = 'b111011000;assign rom[14373] = 'b111011000;assign rom[14374] = 'b111011000;assign rom[14375] = 'b111011000;assign rom[14376] = 'b101111000;assign rom[14377] = 'b000110011;assign rom[14378] = 'b110000010;assign rom[14379] = 'b001101010;assign rom[14380] = 'b001011000;assign rom[14381] = 'b101001000;assign rom[14382] = 'b000101011;assign rom[14383] = 'b110000010;assign rom[14384] = 'b111000000;assign rom[14385] = 'b101001100;assign rom[14386] = 'b001001010;assign rom[14387] = 'b111111000;assign rom[14388] = 'b111101000;assign rom[14389] = 'b101001111;assign rom[14390] = 'b000111010;assign rom[14391] = 'b101110110;assign rom[14392] = 'b101100010;assign rom[14393] = 'b101001100;assign rom[14394] = 'b001001010;assign rom[14395] = 'b111011010;assign rom[14396] = 'b111011010;assign rom[14397] = 'b111011010;assign rom[14398] = 'b111011010;assign rom[14399] = 'b111011000;assign rom[14400] = 'b111011000;assign rom[14401] = 'b111011000;assign rom[14402] = 'b111011000;assign rom[14403] = 'b101111000;assign rom[14404] = 'b000110011;assign rom[14405] = 'b110000010;assign rom[14406] = 'b001101010;assign rom[14407] = 'b001011000;assign rom[14408] = 'b101001000;assign rom[14409] = 'b000101011;assign rom[14410] = 'b110000010;assign rom[14411] = 'b111000000;assign rom[14412] = 'b101001100;assign rom[14413] = 'b001001010;assign rom[14414] = 'b111111000;assign rom[14415] = 'b111101000;assign rom[14416] = 'b101001111;assign rom[14417] = 'b000111010;assign rom[14418] = 'b101110110;assign rom[14419] = 'b101100010;assign rom[14420] = 'b101001100;assign rom[14421] = 'b001001010;assign rom[14422] = 'b111011010;assign rom[14423] = 'b111011010;assign rom[14424] = 'b111011010;assign rom[14425] = 'b111011010;assign rom[14426] = 'b111011000;assign rom[14427] = 'b111011000;assign rom[14428] = 'b111011000;assign rom[14429] = 'b111011000;assign rom[14430] = 'b101111000;assign rom[14431] = 'b000110011;assign rom[14432] = 'b110000010;assign rom[14433] = 'b001101010;assign rom[14434] = 'b001011000;assign rom[14435] = 'b101001000;assign rom[14436] = 'b000101011;assign rom[14437] = 'b110000010;assign rom[14438] = 'b111000000;assign rom[14439] = 'b101001100;assign rom[14440] = 'b001001010;assign rom[14441] = 'b001000110;assign rom[14442] = 'b001100100;assign rom[14443] = 'b101100010;assign rom[14444] = 'b101001100;assign rom[14445] = 'b001001010;assign rom[14446] = 'b111011010;assign rom[14447] = 'b111011010;assign rom[14448] = 'b111011010;assign rom[14449] = 'b111011010;assign rom[14450] = 'b111011000;assign rom[14451] = 'b111011000;assign rom[14452] = 'b111011000;assign rom[14453] = 'b111011000;assign rom[14454] = 'b101111000;assign rom[14455] = 'b000110011;assign rom[14456] = 'b110000010;assign rom[14457] = 'b001101010;assign rom[14458] = 'b001011000;assign rom[14459] = 'b101001000;assign rom[14460] = 'b000101011;assign rom[14461] = 'b110000010;assign rom[14462] = 'b111000000;assign rom[14463] = 'b101001100;assign rom[14464] = 'b001001010;assign rom[14465] = 'b111111000;assign rom[14466] = 'b111101000;assign rom[14467] = 'b101001111;assign rom[14468] = 'b000111010;assign rom[14469] = 'b101110110;assign rom[14470] = 'b101100010;assign rom[14471] = 'b101001100;assign rom[14472] = 'b001001010;assign rom[14473] = 'b111011010;assign rom[14474] = 'b111011010;assign rom[14475] = 'b111011010;assign rom[14476] = 'b111011010;assign rom[14477] = 'b111011000;assign rom[14478] = 'b111011000;assign rom[14479] = 'b111011000;assign rom[14480] = 'b111011000;assign rom[14481] = 'b101111000;assign rom[14482] = 'b000110011;assign rom[14483] = 'b110000010;assign rom[14484] = 'b001101010;assign rom[14485] = 'b001011000;assign rom[14486] = 'b101001000;assign rom[14487] = 'b000101011;assign rom[14488] = 'b110000010;assign rom[14489] = 'b111000000;assign rom[14490] = 'b101001100;assign rom[14491] = 'b001001010;assign rom[14492] = 'b111111000;assign rom[14493] = 'b111101000;assign rom[14494] = 'b101001111;assign rom[14495] = 'b000111010;assign rom[14496] = 'b101110110;assign rom[14497] = 'b101100010;assign rom[14498] = 'b101001100;assign rom[14499] = 'b001001010;assign rom[14500] = 'b111011010;assign rom[14501] = 'b111011010;assign rom[14502] = 'b111011010;assign rom[14503] = 'b111011010;assign rom[14504] = 'b111011000;assign rom[14505] = 'b111011000;assign rom[14506] = 'b111011000;assign rom[14507] = 'b111011000;assign rom[14508] = 'b101111000;assign rom[14509] = 'b000110011;assign rom[14510] = 'b110000010;assign rom[14511] = 'b001101010;assign rom[14512] = 'b001011000;assign rom[14513] = 'b101001000;assign rom[14514] = 'b000101011;assign rom[14515] = 'b110000010;assign rom[14516] = 'b111000000;assign rom[14517] = 'b101001100;assign rom[14518] = 'b001001010;assign rom[14519] = 'b111111000;assign rom[14520] = 'b111101000;assign rom[14521] = 'b101001111;assign rom[14522] = 'b000111010;assign rom[14523] = 'b101110110;assign rom[14524] = 'b101100010;assign rom[14525] = 'b101001100;assign rom[14526] = 'b001001010;assign rom[14527] = 'b111011010;assign rom[14528] = 'b111011010;assign rom[14529] = 'b111011010;assign rom[14530] = 'b111011010;assign rom[14531] = 'b111011000;assign rom[14532] = 'b111011000;assign rom[14533] = 'b111011000;assign rom[14534] = 'b111011000;assign rom[14535] = 'b101111000;assign rom[14536] = 'b000110011;assign rom[14537] = 'b110000010;assign rom[14538] = 'b001101010;assign rom[14539] = 'b001011000;assign rom[14540] = 'b101001000;assign rom[14541] = 'b000101011;assign rom[14542] = 'b110000010;assign rom[14543] = 'b111000000;assign rom[14544] = 'b101001100;assign rom[14545] = 'b001001010;assign rom[14546] = 'b111111000;assign rom[14547] = 'b111101000;assign rom[14548] = 'b101001111;assign rom[14549] = 'b000111010;assign rom[14550] = 'b101110110;assign rom[14551] = 'b101100010;assign rom[14552] = 'b101001100;assign rom[14553] = 'b001001010;assign rom[14554] = 'b111011010;assign rom[14555] = 'b111011010;assign rom[14556] = 'b111011010;assign rom[14557] = 'b111011010;assign rom[14558] = 'b111011000;assign rom[14559] = 'b111011000;assign rom[14560] = 'b111011000;assign rom[14561] = 'b111011000;assign rom[14562] = 'b101111000;assign rom[14563] = 'b000110011;assign rom[14564] = 'b110000010;assign rom[14565] = 'b001101010;assign rom[14566] = 'b001011000;assign rom[14567] = 'b101001000;assign rom[14568] = 'b000101011;assign rom[14569] = 'b110000010;assign rom[14570] = 'b111000000;assign rom[14571] = 'b101001100;assign rom[14572] = 'b001001010;assign rom[14573] = 'b111111000;assign rom[14574] = 'b111101000;assign rom[14575] = 'b101001111;assign rom[14576] = 'b000111010;assign rom[14577] = 'b101110110;assign rom[14578] = 'b101100010;assign rom[14579] = 'b101001100;assign rom[14580] = 'b001001010;assign rom[14581] = 'b111011010;assign rom[14582] = 'b111011010;assign rom[14583] = 'b111011010;assign rom[14584] = 'b111011010;assign rom[14585] = 'b111011000;assign rom[14586] = 'b111011000;assign rom[14587] = 'b111011000;assign rom[14588] = 'b111011000;assign rom[14589] = 'b101111000;assign rom[14590] = 'b000110011;assign rom[14591] = 'b110000010;assign rom[14592] = 'b001101010;assign rom[14593] = 'b001011000;assign rom[14594] = 'b101001000;assign rom[14595] = 'b000101011;assign rom[14596] = 'b110000010;assign rom[14597] = 'b111000000;assign rom[14598] = 'b101001100;assign rom[14599] = 'b001001010;assign rom[14600] = 'b111111000;assign rom[14601] = 'b111101000;assign rom[14602] = 'b101001111;assign rom[14603] = 'b000111010;assign rom[14604] = 'b101110110;assign rom[14605] = 'b101100010;assign rom[14606] = 'b101001100;assign rom[14607] = 'b001001010;assign rom[14608] = 'b111011010;assign rom[14609] = 'b111011010;assign rom[14610] = 'b111011010;assign rom[14611] = 'b111011010;assign rom[14612] = 'b111011000;assign rom[14613] = 'b111011000;assign rom[14614] = 'b111011000;assign rom[14615] = 'b111011000;assign rom[14616] = 'b101111000;assign rom[14617] = 'b000110011;assign rom[14618] = 'b110000010;assign rom[14619] = 'b001101010;assign rom[14620] = 'b001011000;assign rom[14621] = 'b101001000;assign rom[14622] = 'b000101011;assign rom[14623] = 'b110000010;assign rom[14624] = 'b111000000;assign rom[14625] = 'b101001100;assign rom[14626] = 'b001001010;assign rom[14627] = 'b111111000;assign rom[14628] = 'b111101000;assign rom[14629] = 'b101001111;assign rom[14630] = 'b000111010;assign rom[14631] = 'b101110110;assign rom[14632] = 'b101100010;assign rom[14633] = 'b101001100;assign rom[14634] = 'b001001010;assign rom[14635] = 'b111011010;assign rom[14636] = 'b111011010;assign rom[14637] = 'b111011010;assign rom[14638] = 'b111011010;assign rom[14639] = 'b111011000;assign rom[14640] = 'b111011000;assign rom[14641] = 'b111011000;assign rom[14642] = 'b111011000;assign rom[14643] = 'b101111000;assign rom[14644] = 'b000110011;assign rom[14645] = 'b110000010;assign rom[14646] = 'b001101010;assign rom[14647] = 'b001011000;assign rom[14648] = 'b101001000;assign rom[14649] = 'b000101011;assign rom[14650] = 'b110000010;assign rom[14651] = 'b111000000;assign rom[14652] = 'b101001100;assign rom[14653] = 'b001001010;assign rom[14654] = 'b111111000;assign rom[14655] = 'b111101000;assign rom[14656] = 'b101001111;assign rom[14657] = 'b000111010;assign rom[14658] = 'b101110110;assign rom[14659] = 'b101100010;assign rom[14660] = 'b101001100;assign rom[14661] = 'b001001010;assign rom[14662] = 'b111011010;assign rom[14663] = 'b111011010;assign rom[14664] = 'b111011010;assign rom[14665] = 'b111011010;assign rom[14666] = 'b111011000;assign rom[14667] = 'b111011000;assign rom[14668] = 'b111011000;assign rom[14669] = 'b111011000;assign rom[14670] = 'b101111000;assign rom[14671] = 'b000110011;assign rom[14672] = 'b110000010;assign rom[14673] = 'b001101010;assign rom[14674] = 'b001011000;assign rom[14675] = 'b101001000;assign rom[14676] = 'b000101011;assign rom[14677] = 'b110000010;assign rom[14678] = 'b111000000;assign rom[14679] = 'b101001100;assign rom[14680] = 'b001001010;assign rom[14681] = 'b001000110;assign rom[14682] = 'b001100100;assign rom[14683] = 'b101100010;assign rom[14684] = 'b101001100;assign rom[14685] = 'b001001010;assign rom[14686] = 'b111011010;assign rom[14687] = 'b111011010;assign rom[14688] = 'b111011010;assign rom[14689] = 'b111011010;assign rom[14690] = 'b111011000;assign rom[14691] = 'b111011000;assign rom[14692] = 'b111011000;assign rom[14693] = 'b111011000;assign rom[14694] = 'b101111000;assign rom[14695] = 'b000110011;assign rom[14696] = 'b110000010;assign rom[14697] = 'b001101010;assign rom[14698] = 'b001011000;assign rom[14699] = 'b101001000;assign rom[14700] = 'b000101011;assign rom[14701] = 'b110000010;assign rom[14702] = 'b111000000;assign rom[14703] = 'b101001100;assign rom[14704] = 'b001001010;assign rom[14705] = 'b111111000;assign rom[14706] = 'b111101000;assign rom[14707] = 'b101001111;assign rom[14708] = 'b000111010;assign rom[14709] = 'b101110110;assign rom[14710] = 'b101100010;assign rom[14711] = 'b101001100;assign rom[14712] = 'b001001010;assign rom[14713] = 'b111011010;assign rom[14714] = 'b111011010;assign rom[14715] = 'b111011010;assign rom[14716] = 'b111011010;assign rom[14717] = 'b111011000;assign rom[14718] = 'b111011000;assign rom[14719] = 'b111011000;assign rom[14720] = 'b111011000;assign rom[14721] = 'b101111000;assign rom[14722] = 'b000110011;assign rom[14723] = 'b110000010;assign rom[14724] = 'b001101010;assign rom[14725] = 'b001011000;assign rom[14726] = 'b101001000;assign rom[14727] = 'b000101011;assign rom[14728] = 'b110000010;assign rom[14729] = 'b111000000;assign rom[14730] = 'b101001100;assign rom[14731] = 'b001001010;assign rom[14732] = 'b111111000;assign rom[14733] = 'b111101000;assign rom[14734] = 'b101001111;assign rom[14735] = 'b000111010;assign rom[14736] = 'b101110110;assign rom[14737] = 'b101100010;assign rom[14738] = 'b101001100;assign rom[14739] = 'b001001010;assign rom[14740] = 'b111011010;assign rom[14741] = 'b111011010;assign rom[14742] = 'b111011010;assign rom[14743] = 'b111011010;assign rom[14744] = 'b111011000;assign rom[14745] = 'b111011000;assign rom[14746] = 'b111011000;assign rom[14747] = 'b111011000;assign rom[14748] = 'b101111000;assign rom[14749] = 'b000110011;assign rom[14750] = 'b110000010;assign rom[14751] = 'b001101010;assign rom[14752] = 'b001011000;assign rom[14753] = 'b101001000;assign rom[14754] = 'b000101011;assign rom[14755] = 'b110000010;assign rom[14756] = 'b111000000;assign rom[14757] = 'b101001100;assign rom[14758] = 'b001001010;assign rom[14759] = 'b111111000;assign rom[14760] = 'b111101000;assign rom[14761] = 'b101001111;assign rom[14762] = 'b000111010;assign rom[14763] = 'b101110110;assign rom[14764] = 'b101100010;assign rom[14765] = 'b101001100;assign rom[14766] = 'b001001010;assign rom[14767] = 'b111011010;assign rom[14768] = 'b111011010;assign rom[14769] = 'b111011010;assign rom[14770] = 'b111011010;assign rom[14771] = 'b111011000;assign rom[14772] = 'b111011000;assign rom[14773] = 'b111011000;assign rom[14774] = 'b111011000;assign rom[14775] = 'b101111000;assign rom[14776] = 'b000110011;assign rom[14777] = 'b110000010;assign rom[14778] = 'b001101010;assign rom[14779] = 'b001011000;assign rom[14780] = 'b101001000;assign rom[14781] = 'b000101011;assign rom[14782] = 'b110000010;assign rom[14783] = 'b111000000;assign rom[14784] = 'b101001100;assign rom[14785] = 'b001001010;assign rom[14786] = 'b111111000;assign rom[14787] = 'b111101000;assign rom[14788] = 'b101001111;assign rom[14789] = 'b000111010;assign rom[14790] = 'b101110110;assign rom[14791] = 'b101100010;assign rom[14792] = 'b101001100;assign rom[14793] = 'b001001010;assign rom[14794] = 'b111011010;assign rom[14795] = 'b111011010;assign rom[14796] = 'b111011010;assign rom[14797] = 'b111011010;assign rom[14798] = 'b111011000;assign rom[14799] = 'b111011000;assign rom[14800] = 'b111011000;assign rom[14801] = 'b111011000;assign rom[14802] = 'b101111000;assign rom[14803] = 'b000110011;assign rom[14804] = 'b110000010;assign rom[14805] = 'b001101010;assign rom[14806] = 'b001011000;assign rom[14807] = 'b101001000;assign rom[14808] = 'b000101011;assign rom[14809] = 'b110000010;assign rom[14810] = 'b111000000;assign rom[14811] = 'b101001100;assign rom[14812] = 'b001001010;assign rom[14813] = 'b111111000;assign rom[14814] = 'b111101000;assign rom[14815] = 'b101001111;assign rom[14816] = 'b000111010;assign rom[14817] = 'b101110110;assign rom[14818] = 'b101100010;assign rom[14819] = 'b101001100;assign rom[14820] = 'b001001010;assign rom[14821] = 'b111011010;assign rom[14822] = 'b111011010;assign rom[14823] = 'b111011010;assign rom[14824] = 'b111011010;assign rom[14825] = 'b111011000;assign rom[14826] = 'b111011000;assign rom[14827] = 'b111011000;assign rom[14828] = 'b111011000;assign rom[14829] = 'b101111000;assign rom[14830] = 'b000110011;assign rom[14831] = 'b110000010;assign rom[14832] = 'b001101010;assign rom[14833] = 'b001011000;assign rom[14834] = 'b101001000;assign rom[14835] = 'b000101011;assign rom[14836] = 'b110000010;assign rom[14837] = 'b111000000;assign rom[14838] = 'b101001100;assign rom[14839] = 'b001001010;assign rom[14840] = 'b111111000;assign rom[14841] = 'b111101000;assign rom[14842] = 'b101001111;assign rom[14843] = 'b000111010;assign rom[14844] = 'b101110110;assign rom[14845] = 'b101100010;assign rom[14846] = 'b101001100;assign rom[14847] = 'b001001010;assign rom[14848] = 'b111011010;assign rom[14849] = 'b111011010;assign rom[14850] = 'b111011010;assign rom[14851] = 'b111011010;assign rom[14852] = 'b111011000;assign rom[14853] = 'b111011000;assign rom[14854] = 'b111011000;assign rom[14855] = 'b111011000;assign rom[14856] = 'b101111000;assign rom[14857] = 'b000110011;assign rom[14858] = 'b110000010;assign rom[14859] = 'b001101010;assign rom[14860] = 'b001011000;assign rom[14861] = 'b101001000;assign rom[14862] = 'b000101011;assign rom[14863] = 'b110000010;assign rom[14864] = 'b111000000;assign rom[14865] = 'b101001100;assign rom[14866] = 'b001001010;assign rom[14867] = 'b111111000;assign rom[14868] = 'b111101000;assign rom[14869] = 'b101001111;assign rom[14870] = 'b000111010;assign rom[14871] = 'b101110110;assign rom[14872] = 'b101100010;assign rom[14873] = 'b101001100;assign rom[14874] = 'b001001010;assign rom[14875] = 'b111011010;assign rom[14876] = 'b111011010;assign rom[14877] = 'b111011010;assign rom[14878] = 'b111011010;assign rom[14879] = 'b111011000;assign rom[14880] = 'b111011000;assign rom[14881] = 'b111011000;assign rom[14882] = 'b111011000;assign rom[14883] = 'b101111000;assign rom[14884] = 'b000110011;assign rom[14885] = 'b110000010;assign rom[14886] = 'b001101010;assign rom[14887] = 'b001011000;assign rom[14888] = 'b101001000;assign rom[14889] = 'b000101011;assign rom[14890] = 'b110000010;assign rom[14891] = 'b111000000;assign rom[14892] = 'b101001100;assign rom[14893] = 'b001001010;assign rom[14894] = 'b111111000;assign rom[14895] = 'b111101000;assign rom[14896] = 'b101001111;assign rom[14897] = 'b000111010;assign rom[14898] = 'b101110110;assign rom[14899] = 'b101100010;assign rom[14900] = 'b101001100;assign rom[14901] = 'b001001010;assign rom[14902] = 'b111011010;assign rom[14903] = 'b111011010;assign rom[14904] = 'b111011010;assign rom[14905] = 'b111011010;assign rom[14906] = 'b111011000;assign rom[14907] = 'b111011000;assign rom[14908] = 'b111011000;assign rom[14909] = 'b111011000;assign rom[14910] = 'b101111000;assign rom[14911] = 'b000110011;assign rom[14912] = 'b110000010;assign rom[14913] = 'b001101010;assign rom[14914] = 'b001011000;assign rom[14915] = 'b101001000;assign rom[14916] = 'b000101011;assign rom[14917] = 'b110000010;assign rom[14918] = 'b111000000;assign rom[14919] = 'b101001100;assign rom[14920] = 'b001001010;assign rom[14921] = 'b001000110;assign rom[14922] = 'b001100100;assign rom[14923] = 'b101100010;assign rom[14924] = 'b101001100;assign rom[14925] = 'b001001010;assign rom[14926] = 'b111011010;assign rom[14927] = 'b111011010;assign rom[14928] = 'b111011010;assign rom[14929] = 'b111011010;assign rom[14930] = 'b111011000;assign rom[14931] = 'b111011000;assign rom[14932] = 'b111011000;assign rom[14933] = 'b111011000;assign rom[14934] = 'b101111000;assign rom[14935] = 'b000110011;assign rom[14936] = 'b110000010;assign rom[14937] = 'b001101010;assign rom[14938] = 'b001011000;assign rom[14939] = 'b101001000;assign rom[14940] = 'b000101011;assign rom[14941] = 'b110000010;assign rom[14942] = 'b111000000;assign rom[14943] = 'b101001100;assign rom[14944] = 'b001001010;assign rom[14945] = 'b111111000;assign rom[14946] = 'b111101000;assign rom[14947] = 'b101001111;assign rom[14948] = 'b000111010;assign rom[14949] = 'b101110110;assign rom[14950] = 'b101100010;assign rom[14951] = 'b101001100;assign rom[14952] = 'b001001010;assign rom[14953] = 'b111011010;assign rom[14954] = 'b111011010;assign rom[14955] = 'b111011010;assign rom[14956] = 'b111011010;assign rom[14957] = 'b111011000;assign rom[14958] = 'b111011000;assign rom[14959] = 'b111011000;assign rom[14960] = 'b111011000;assign rom[14961] = 'b101111000;assign rom[14962] = 'b000110011;assign rom[14963] = 'b110000010;assign rom[14964] = 'b001101010;assign rom[14965] = 'b001011000;assign rom[14966] = 'b101001000;assign rom[14967] = 'b000101011;assign rom[14968] = 'b110000010;assign rom[14969] = 'b111000000;assign rom[14970] = 'b101001100;assign rom[14971] = 'b001001010;assign rom[14972] = 'b111111000;assign rom[14973] = 'b111101000;assign rom[14974] = 'b101001111;assign rom[14975] = 'b000111010;assign rom[14976] = 'b101110110;assign rom[14977] = 'b101100010;assign rom[14978] = 'b101001100;assign rom[14979] = 'b001001010;assign rom[14980] = 'b111011010;assign rom[14981] = 'b111011010;assign rom[14982] = 'b111011010;assign rom[14983] = 'b111011010;assign rom[14984] = 'b111011000;assign rom[14985] = 'b111011000;assign rom[14986] = 'b111011000;assign rom[14987] = 'b111011000;assign rom[14988] = 'b101111000;assign rom[14989] = 'b000110011;assign rom[14990] = 'b110000010;assign rom[14991] = 'b001101010;assign rom[14992] = 'b001011000;assign rom[14993] = 'b101001000;assign rom[14994] = 'b000101011;assign rom[14995] = 'b110000010;assign rom[14996] = 'b111000000;assign rom[14997] = 'b101001100;assign rom[14998] = 'b001001010;assign rom[14999] = 'b111111000;assign rom[15000] = 'b111101000;assign rom[15001] = 'b101001111;assign rom[15002] = 'b000111010;assign rom[15003] = 'b101110110;assign rom[15004] = 'b101100010;assign rom[15005] = 'b101001100;assign rom[15006] = 'b001001010;assign rom[15007] = 'b111011010;assign rom[15008] = 'b111011010;assign rom[15009] = 'b111011010;assign rom[15010] = 'b111011010;assign rom[15011] = 'b111011000;assign rom[15012] = 'b111011000;assign rom[15013] = 'b111011000;assign rom[15014] = 'b111011000;assign rom[15015] = 'b101111000;assign rom[15016] = 'b000110011;assign rom[15017] = 'b110000010;assign rom[15018] = 'b001101010;assign rom[15019] = 'b001011000;assign rom[15020] = 'b101001000;assign rom[15021] = 'b000101011;assign rom[15022] = 'b110000010;assign rom[15023] = 'b111000000;assign rom[15024] = 'b101001100;assign rom[15025] = 'b001001010;assign rom[15026] = 'b111111000;assign rom[15027] = 'b111101000;assign rom[15028] = 'b101001111;assign rom[15029] = 'b000111010;assign rom[15030] = 'b101110110;assign rom[15031] = 'b101100010;assign rom[15032] = 'b101001100;assign rom[15033] = 'b001001010;assign rom[15034] = 'b111011010;assign rom[15035] = 'b111011010;assign rom[15036] = 'b111011010;assign rom[15037] = 'b111011010;assign rom[15038] = 'b111011000;assign rom[15039] = 'b111011000;assign rom[15040] = 'b111011000;assign rom[15041] = 'b111011000;assign rom[15042] = 'b101111000;assign rom[15043] = 'b000110011;assign rom[15044] = 'b110000010;assign rom[15045] = 'b001101010;assign rom[15046] = 'b001011000;assign rom[15047] = 'b101001000;assign rom[15048] = 'b000101011;assign rom[15049] = 'b110000010;assign rom[15050] = 'b111000000;assign rom[15051] = 'b101001100;assign rom[15052] = 'b001001010;assign rom[15053] = 'b111111000;assign rom[15054] = 'b111101000;assign rom[15055] = 'b101001111;assign rom[15056] = 'b000111010;assign rom[15057] = 'b101110110;assign rom[15058] = 'b101100010;assign rom[15059] = 'b101001100;assign rom[15060] = 'b001001010;assign rom[15061] = 'b111011010;assign rom[15062] = 'b111011010;assign rom[15063] = 'b111011010;assign rom[15064] = 'b111011010;assign rom[15065] = 'b111011000;assign rom[15066] = 'b111011000;assign rom[15067] = 'b111011000;assign rom[15068] = 'b111011000;assign rom[15069] = 'b101111000;assign rom[15070] = 'b000110011;assign rom[15071] = 'b110000010;assign rom[15072] = 'b001101010;assign rom[15073] = 'b001011000;assign rom[15074] = 'b101001000;assign rom[15075] = 'b000101011;assign rom[15076] = 'b110000010;assign rom[15077] = 'b111000000;assign rom[15078] = 'b101001100;assign rom[15079] = 'b001001010;assign rom[15080] = 'b111111000;assign rom[15081] = 'b111101000;assign rom[15082] = 'b101001111;assign rom[15083] = 'b000111010;assign rom[15084] = 'b101110110;assign rom[15085] = 'b101100010;assign rom[15086] = 'b101001100;assign rom[15087] = 'b001001010;assign rom[15088] = 'b111011010;assign rom[15089] = 'b111011010;assign rom[15090] = 'b111011010;assign rom[15091] = 'b111011010;assign rom[15092] = 'b111011000;assign rom[15093] = 'b111011000;assign rom[15094] = 'b111011000;assign rom[15095] = 'b111011000;assign rom[15096] = 'b101111000;assign rom[15097] = 'b000110011;assign rom[15098] = 'b110000010;assign rom[15099] = 'b001101010;assign rom[15100] = 'b001011000;assign rom[15101] = 'b101001000;assign rom[15102] = 'b000101011;assign rom[15103] = 'b110000010;assign rom[15104] = 'b111000000;assign rom[15105] = 'b101001100;assign rom[15106] = 'b001001010;assign rom[15107] = 'b111111000;assign rom[15108] = 'b111101000;assign rom[15109] = 'b101001111;assign rom[15110] = 'b000111010;assign rom[15111] = 'b101110110;assign rom[15112] = 'b101100010;assign rom[15113] = 'b101001100;assign rom[15114] = 'b001001010;assign rom[15115] = 'b111011010;assign rom[15116] = 'b111011010;assign rom[15117] = 'b111011010;assign rom[15118] = 'b111011010;assign rom[15119] = 'b111011000;assign rom[15120] = 'b111011000;assign rom[15121] = 'b111011000;assign rom[15122] = 'b111011000;assign rom[15123] = 'b101111000;assign rom[15124] = 'b000110011;assign rom[15125] = 'b110000010;assign rom[15126] = 'b001101010;assign rom[15127] = 'b001011000;assign rom[15128] = 'b101001000;assign rom[15129] = 'b000101011;assign rom[15130] = 'b110000010;assign rom[15131] = 'b111000000;assign rom[15132] = 'b101001100;assign rom[15133] = 'b001001010;assign rom[15134] = 'b111111000;assign rom[15135] = 'b111101000;assign rom[15136] = 'b101001111;assign rom[15137] = 'b000111010;assign rom[15138] = 'b101110110;assign rom[15139] = 'b101100010;assign rom[15140] = 'b101001100;assign rom[15141] = 'b001001010;assign rom[15142] = 'b111011010;assign rom[15143] = 'b111011010;assign rom[15144] = 'b111011010;assign rom[15145] = 'b111011010;assign rom[15146] = 'b111011000;assign rom[15147] = 'b111011000;assign rom[15148] = 'b111011000;assign rom[15149] = 'b111011000;assign rom[15150] = 'b101111000;assign rom[15151] = 'b000110011;assign rom[15152] = 'b110000010;assign rom[15153] = 'b001101010;assign rom[15154] = 'b001011000;assign rom[15155] = 'b101001000;assign rom[15156] = 'b000101011;assign rom[15157] = 'b110000010;assign rom[15158] = 'b111000000;assign rom[15159] = 'b101001100;assign rom[15160] = 'b001001010;assign rom[15161] = 'b001000110;assign rom[15162] = 'b001100100;
endmodule
