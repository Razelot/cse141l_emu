`timescale 1ns / 1ps

module reg_file #(parameter num_regs = 12, reg_width = 8)
(
  input clk,
  input read, write, write_car,
  input [$clog2(num_regs)-1:0] rt_addr, rs_addr, rd_addr,
  input [reg_width-1:0] rd_in, car_in
  output logic [reg_width-1:0] rt_out, rs_out);

  // register array
  logic [reg_width-1:0] regs [num_regs-1:0];

  logic allow_write;

  // cannot write reg[0]
  assign allow_write = rd_addr != 8'b0000 && write;

  always_ff @ (posedge clk ) begin

    if(read) begin
    rt_out <= regs[rt_addr];
    rs_out <= regs[rs_addr];
    end

    if(allow_write)
    regs[rd_addr] <= rd_in;

    if(write_car)
    regs[11] <= car_in;

  end

  endmodule
